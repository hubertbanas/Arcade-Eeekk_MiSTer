library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_0 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"01",X"53",X"A3",X"BF",X"B5",X"A3",X"3D",X"B5",X"10",X"9F",X"0E",X"A1",X"D7",X"37",X"88",X"E9",
		X"AF",X"10",X"F9",X"5C",X"64",X"BB",X"10",X"FF",X"98",X"7D",X"D2",X"07",X"37",X"7D",X"17",X"77",
		X"37",X"40",X"03",X"36",X"EC",X"22",X"B5",X"34",X"5F",X"27",X"E0",X"98",X"13",X"98",X"5D",X"53",
		X"A3",X"9B",X"B5",X"E6",X"19",X"03",X"9F",X"F8",X"45",X"5D",X"55",X"4D",X"A2",X"C2",X"FC",X"4B",
		X"38",X"08",X"BF",X"10",X"FB",X"54",X"B2",X"09",X"55",X"33",X"34",X"57",X"E1",X"29",X"98",X"41",
		X"A2",X"41",X"C7",X"DB",X"DB",X"45",X"A2",X"0A",X"FC",X"4B",X"AE",X"AB",X"A2",X"6E",X"FC",X"4B",
		X"AE",X"F6",X"E0",X"C6",X"18",X"F8",X"AF",X"BB",X"79",X"FF",X"5C",X"44",X"BF",X"E2",X"69",X"73",
		X"79",X"EB",X"BB",X"9B",X"8B",X"E0",X"71",X"B6",X"71",X"24",X"4C",X"FD",X"B6",X"9E",X"E0",X"5C",
		X"44",X"BF",X"E0",X"BB",X"9B",X"8B",X"E0",X"BB",X"9B",X"8B",X"05",X"C6",X"AF",X"59",X"A2",X"2A",
		X"FC",X"4B",X"AF",X"87",X"A2",X"0F",X"F8",X"4B",X"AE",X"8A",X"D9",X"8F",X"BA",X"D8",X"8B",X"8B",
		X"F0",X"8B",X"F1",X"8B",X"E0",X"69",X"DA",X"8B",X"5D",X"4D",X"55",X"C6",X"D0",X"DB",X"DB",X"1B",
		X"DB",X"DB",X"F3",X"BF",X"D0",X"8F",X"BA",X"8A",X"96",X"15",X"08",X"9F",X"BB",X"DF",X"5C",X"52",
		X"FF",X"0D",X"1D",X"B7",X"14",X"8F",X"DB",X"FC",X"C7",X"8B",X"E3",X"BF",X"8B",X"C7",X"AF",X"9B",
		X"5C",X"80",X"C2",X"5C",X"F7",X"BE",X"5C",X"E3",X"9F",X"10",X"9F",X"1F",X"15",X"1D",X"41",X"F3",
		X"FD",X"B5",X"E6",X"F3",X"FD",X"B5",X"10",X"FD",X"05",X"00",X"1C",X"A2",X"2A",X"FC",X"4B",X"AF",
		X"75",X"8F",X"21",X"D8",X"53",X"FB",X"FE",X"C1",X"8B",X"B7",X"64",X"B6",X"3C",X"5D",X"D9",X"60",
		X"FD",X"A6",X"93",X"A2",X"2D",X"DC",X"60",X"9B",X"FA",X"A4",X"AE",X"BE",X"60",X"BB",X"FA",X"BF",
		X"AE",X"BB",X"FA",X"E6",X"A4",X"1F",X"1D",X"B3",X"93",X"8B",X"E0",X"B3",X"93",X"8B",X"1C",X"45",
		X"5D",X"FB",X"40",X"A2",X"DE",X"FC",X"18",X"C1",X"AF",X"BB",X"FB",X"42",X"5C",X"96",X"BB",X"2F",
		X"A3",X"DE",X"FC",X"1D",X"05",X"1C",X"45",X"4D",X"A2",X"4A",X"FC",X"4B",X"AF",X"96",X"5C",X"B0",
		X"9F",X"A2",X"BF",X"B5",X"69",X"B7",X"38",X"91",X"97",X"A2",X"0A",X"FC",X"4B",X"AF",X"BE",X"A2",
		X"BD",X"B5",X"69",X"B7",X"38",X"91",X"97",X"0D",X"05",X"1C",X"A2",X"DA",X"FC",X"4B",X"AE",X"EE",
		X"A2",X"BF",X"B5",X"18",X"C8",X"3D",X"53",X"A3",X"DA",X"FC",X"E6",X"A3",X"97",X"FC",X"5C",X"63",
		X"DB",X"E2",X"BF",X"5C",X"A6",X"BA",X"8F",X"A2",X"FC",X"E0",X"60",X"16",X"3C",X"79",X"9F",X"CB",
		X"C1",X"E2",X"DA",X"A3",X"FE",X"FC",X"E2",X"9F",X"A3",X"DB",X"B5",X"1C",X"8F",X"FE",X"FC",X"C7",
		X"3D",X"E3",X"9F",X"A2",X"BF",X"B5",X"18",X"C8",X"3C",X"53",X"A3",X"DB",X"B5",X"E6",X"A3",X"DA",
		X"FC",X"1C",X"5C",X"79",X"9E",X"5C",X"63",X"DB",X"E2",X"BE",X"5C",X"A6",X"BA",X"5C",X"A6",X"9B",
		X"19",X"BB",X"82",X"A3",X"16",X"FC",X"A3",X"4F",X"F8",X"A3",X"DA",X"FC",X"A3",X"B3",X"FC",X"8F",
		X"F8",X"FC",X"E3",X"91",X"8B",X"E3",X"9C",X"8B",X"E3",X"FD",X"8B",X"E3",X"BF",X"8B",X"E3",X"9F",
		X"8B",X"E3",X"BF",X"A2",X"BD",X"B5",X"18",X"C0",X"E2",X"9F",X"AE",X"9F",X"53",X"A3",X"0A",X"FC",
		X"19",X"28",X"C2",X"45",X"69",X"25",X"DA",X"DA",X"DA",X"DA",X"D9",X"05",X"69",X"DA",X"D8",X"1C",
		X"45",X"A2",X"37",X"FC",X"B6",X"FF",X"45",X"A2",X"FF",X"DC",X"5D",X"D9",X"A2",X"0A",X"FC",X"4B",
		X"AE",X"DA",X"A4",X"FB",X"BF",X"60",X"9F",X"AE",X"9F",X"FF",X"A4",X"A3",X"9B",X"B5",X"A3",X"6E",
		X"FC",X"1D",X"05",X"1C",X"A2",X"37",X"FC",X"B6",X"9B",X"A2",X"FF",X"DC",X"5D",X"D9",X"A2",X"0A",
		X"FC",X"4B",X"AE",X"92",X"A4",X"60",X"9F",X"AE",X"F3",X"A2",X"BD",X"B5",X"D9",X"69",X"DA",X"D8",
		X"A4",X"69",X"B7",X"DB",X"07",X"D8",X"A2",X"BF",X"B5",X"69",X"3F",X"DA",X"07",X"1D",X"1C",X"A2",
		X"BF",X"B5",X"69",X"DA",X"D8",X"A2",X"BD",X"B5",X"69",X"AD",X"B6",X"25",X"5C",X"D5",X"BB",X"FB",
		X"F2",X"5C",X"9E",X"9B",X"1C",X"5C",X"8C",X"BB",X"5C",X"A0",X"BB",X"5C",X"4E",X"BB",X"1C",X"5C",
		X"1A",X"BB",X"5C",X"76",X"BB",X"5C",X"23",X"BB",X"1C",X"8F",X"39",X"99",X"9F",X"9F",X"F6",X"5C",
		X"26",X"BB",X"8F",X"29",X"99",X"9F",X"9F",X"F6",X"B6",X"E2",X"8F",X"BB",X"BD",X"9F",X"9F",X"F6",
		X"5C",X"26",X"BB",X"8F",X"AB",X"BD",X"9F",X"9F",X"F6",X"B6",X"CE",X"8F",X"39",X"D9",X"9F",X"9F",
		X"F6",X"5C",X"26",X"BB",X"8F",X"29",X"D9",X"9F",X"9F",X"F6",X"B6",X"F6",X"8F",X"BB",X"FD",X"9F",
		X"9F",X"F6",X"5C",X"26",X"BB",X"8F",X"AB",X"FD",X"9F",X"9F",X"F6",X"B6",X"9A",X"8F",X"BD",X"BD",
		X"B6",X"9B",X"8F",X"BD",X"FD",X"9F",X"FF",X"3F",X"C1",X"8B",X"B7",X"64",X"A3",X"3D",X"B5",X"DE",
		X"AF",X"61",X"1C",X"FB",X"E6",X"5C",X"0D",X"BB",X"E2",X"9F",X"A3",X"BF",X"B5",X"00",X"A2",X"BE",
		X"FC",X"4B",X"AF",X"05",X"A3",X"3D",X"B5",X"E6",X"A3",X"BE",X"FC",X"B7",X"2C",X"DE",X"AF",X"09",
		X"1C",X"45",X"A2",X"A2",X"FC",X"4B",X"AF",X"BB",X"05",X"1C",X"87",X"25",X"D8",X"53",X"A3",X"B7",
		X"FC",X"A3",X"C2",X"FC",X"E6",X"A3",X"BF",X"B5",X"00",X"19",X"F5",X"B2",X"5D",X"FA",X"BF",X"DE",
		X"AF",X"44",X"A3",X"3D",X"B5",X"B7",X"24",X"1D",X"1C",X"45",X"5D",X"A4",X"A3",X"DB",X"FC",X"E2",
		X"9F",X"A3",X"BF",X"B5",X"00",X"A3",X"3D",X"B5",X"A2",X"DB",X"FC",X"4B",X"AF",X"05",X"1D",X"05",
		X"1C",X"45",X"E2",X"9F",X"A3",X"BE",X"FC",X"E2",X"9F",X"A3",X"BF",X"B5",X"00",X"A3",X"3D",X"B5",
		X"A2",X"BE",X"FC",X"4B",X"AF",X"05",X"05",X"1C",X"4D",X"8F",X"BC",X"9B",X"5F",X"C8",X"E2",X"BF",
		X"7F",X"C9",X"F9",X"5C",X"9E",X"9B",X"0D",X"1C",X"9F",X"40",X"40",X"A1",X"6A",X"34",X"E6",X"F5",
		X"40",X"74",X"4D",X"8F",X"BC",X"9B",X"5F",X"C8",X"E2",X"BF",X"7E",X"C9",X"F8",X"18",X"86",X"8F",
		X"38",X"F8",X"5C",X"CC",X"9B",X"5C",X"CC",X"9B",X"DE",X"AF",X"65",X"0D",X"1C",X"FB",X"9B",X"5D",
		X"A4",X"4C",X"FD",X"79",X"FB",X"A3",X"C6",X"D8",X"4D",X"F9",X"8B",X"F8",X"8B",X"8B",X"5C",X"B9",
		X"AB",X"0D",X"97",X"9A",X"BF",X"96",X"1D",X"B7",X"69",X"5C",X"8F",X"9B",X"1C",X"55",X"E2",X"9F",
		X"A3",X"FB",X"FC",X"B2",X"5C",X"4B",X"9B",X"93",X"B2",X"5C",X"4B",X"9B",X"93",X"53",X"A3",X"FB",
		X"FC",X"B2",X"5C",X"4B",X"9B",X"15",X"1C",X"5D",X"5C",X"09",X"9F",X"A4",X"5C",X"47",X"9B",X"84",
		X"5C",X"47",X"9B",X"1D",X"1C",X"55",X"D0",X"A2",X"FB",X"FC",X"D1",X"4B",X"AE",X"9E",X"80",X"4B",
		X"E2",X"BF",X"AF",X"9B",X"F2",X"35",X"A0",X"A3",X"FB",X"FC",X"80",X"79",X"A7",X"15",X"55",X"C1",
		X"4D",X"97",X"BF",X"FF",X"96",X"A2",X"BF",X"FC",X"C1",X"0D",X"A2",X"4F",X"F8",X"4B",X"97",X"40",
		X"40",X"AE",X"9B",X"97",X"2D",X"40",X"96",X"15",X"1C",X"5D",X"55",X"5C",X"09",X"9F",X"A4",X"60",
		X"BA",X"F3",X"A7",X"A6",X"BB",X"F3",X"C3",X"3B",X"5C",X"78",X"9B",X"84",X"60",X"BA",X"F3",X"A7",
		X"A6",X"BB",X"F3",X"C3",X"3B",X"5C",X"78",X"9B",X"15",X"1D",X"1C",X"84",X"C0",X"08",X"10",X"2A",
		X"87",X"63",X"75",X"0B",X"5C",X"9B",X"97",X"53",X"74",X"86",X"C0",X"72",X"F7",X"29",X"72",X"FF",
		X"2D",X"72",X"B5",X"34",X"6E",X"72",X"35",X"2D",X"72",X"15",X"2D",X"4D",X"77",X"97",X"94",X"5C",
		X"2E",X"A3",X"4A",X"03",X"9F",X"C1",X"96",X"B7",X"64",X"1C",X"45",X"F8",X"1F",X"C1",X"05",X"96",
		X"B7",X"24",X"1C",X"5D",X"9F",X"9F",X"BF",X"B6",X"FF",X"5D",X"9F",X"2D",X"40",X"4C",X"99",X"BB",
		X"FC",X"45",X"AB",X"FF",X"FC",X"5D",X"FA",X"A3",X"01",X"4C",X"BD",X"78",X"4D",X"8F",X"35",X"00",
		X"1D",X"60",X"40",X"AE",X"D7",X"C1",X"5D",X"4D",X"9F",X"BF",X"FF",X"9E",X"A2",X"BF",X"FC",X"C1",
		X"0D",X"1D",X"93",X"4C",X"98",X"BB",X"FC",X"9E",X"B6",X"10",X"93",X"FA",X"F7",X"01",X"4C",X"BD",
		X"78",X"6D",X"50",X"8F",X"35",X"00",X"60",X"40",X"AF",X"9B",X"05",X"1D",X"1C",X"60",X"60",X"AF",
		X"9E",X"AA",X"FF",X"FC",X"8B",X"AB",X"FF",X"FC",X"B6",X"02",X"A3",X"BF",X"FC",X"B6",X"63",X"A4",
		X"BE",X"B6",X"DB",X"F9",X"A4",X"BE",X"8B",X"F8",X"8B",X"08",X"B2",X"93",X"60",X"AF",X"AE",X"9F",
		X"C1",X"5D",X"4D",X"9F",X"BF",X"FF",X"9E",X"B2",X"93",X"4B",X"AE",X"9F",X"C1",X"0D",X"8A",X"1D",
		X"B7",X"2C",X"BE",X"D9",X"BE",X"5D",X"E2",X"2D",X"3F",X"FB",X"40",X"D8",X"9E",X"1D",X"DE",X"AF",
		X"14",X"1C",X"4D",X"01",X"97",X"0D",X"ED",X"9F",X"FF",X"9E",X"4C",X"AC",X"57",X"90",X"65",X"98",
		X"27",X"91",X"55",X"4F",X"4D",X"97",X"9B",X"DF",X"8F",X"32",X"B9",X"5C",X"9C",X"FF",X"A2",X"9F",
		X"FC",X"A3",X"BF",X"FC",X"53",X"A3",X"FB",X"FC",X"A2",X"A2",X"FC",X"8F",X"22",X"9D",X"5C",X"4B",
		X"9B",X"0D",X"1C",X"8A",X"45",X"11",X"30",X"05",X"25",X"1D",X"24",X"8A",X"8A",X"A2",X"FF",X"DC",
		X"60",X"9F",X"AF",X"BE",X"8F",X"44",X"99",X"97",X"56",X"FC",X"B6",X"FB",X"8F",X"49",X"99",X"97",
		X"2F",X"FC",X"53",X"A3",X"4F",X"F8",X"5C",X"5E",X"9B",X"E2",X"9F",X"A3",X"4F",X"F8",X"1C",X"45",
		X"55",X"4D",X"45",X"A2",X"B7",X"FC",X"60",X"9F",X"38",X"ED",X"DF",X"97",X"52",X"FC",X"8F",X"4B",
		X"FC",X"A2",X"FF",X"DC",X"60",X"9F",X"AE",X"FB",X"97",X"2B",X"FC",X"8F",X"0E",X"FC",X"05",X"4D",
		X"C8",X"B2",X"1F",X"CB",X"B3",X"92",X"B2",X"3E",X"CB",X"B3",X"92",X"B2",X"5E",X"CB",X"B3",X"0D",
		X"5C",X"8C",X"DF",X"45",X"05",X"0D",X"15",X"05",X"1C",X"A2",X"36",X"FC",X"D8",X"B2",X"06",X"34",
		X"E0",X"4B",X"3C",X"8A",X"E7",X"5C",X"1F",X"DF",X"E2",X"F7",X"5C",X"A6",X"BA",X"8B",X"E3",X"BF",
		X"1C",X"A2",X"FF",X"DC",X"60",X"9F",X"AF",X"FE",X"4D",X"9F",X"6B",X"FC",X"97",X"50",X"40",X"8F",
		X"D6",X"BD",X"B6",X"BA",X"4D",X"9F",X"2E",X"FC",X"97",X"0D",X"40",X"8F",X"BB",X"BD",X"A2",X"4A",
		X"FC",X"4B",X"AF",X"EB",X"BA",X"4B",X"AE",X"AB",X"60",X"9E",X"A6",X"BB",X"E2",X"BE",X"D9",X"E3",
		X"9F",X"55",X"97",X"AF",X"BF",X"96",X"E2",X"9E",X"C1",X"4D",X"97",X"BF",X"FF",X"96",X"E6",X"C1",
		X"97",X"2D",X"40",X"96",X"C1",X"0D",X"15",X"96",X"B7",X"4D",X"0D",X"1C",X"A2",X"FF",X"DC",X"60",
		X"9F",X"AF",X"9A",X"8F",X"0F",X"99",X"97",X"3B",X"99",X"9F",X"DB",X"DC",X"B6",X"9E",X"8F",X"1D",
		X"BD",X"97",X"3B",X"BD",X"9F",X"BA",X"DC",X"55",X"97",X"65",X"DF",X"5C",X"9C",X"FF",X"0D",X"BA",
		X"5C",X"4B",X"9B",X"1C",X"2D",X"05",X"20",X"05",X"2D",X"8A",X"8A",X"55",X"4D",X"97",X"9E",X"FB",
		X"8F",X"A9",X"B9",X"5C",X"9C",X"FF",X"0D",X"15",X"1C",X"8A",X"58",X"65",X"45",X"45",X"45",X"45",
		X"45",X"45",X"41",X"8A",X"AA",X"61",X"8A",X"51",X"05",X"05",X"05",X"19",X"19",X"57",X"8A",X"58",
		X"69",X"8A",X"AA",X"6D",X"4D",X"4D",X"4D",X"4D",X"4D",X"4D",X"49",X"8A",X"8A",X"45",X"01",X"10",
		X"49",X"0D",X"05",X"0F",X"41",X"DF",X"69",X"A8",X"E9",X"F4",X"83",X"DB",X"F5",X"26",X"E6",X"F3",
		X"C2",X"AC",X"F3",X"7A",X"AC",X"10",X"F3",X"00",X"8F",X"7B",X"F8",X"E3",X"FB",X"8B",X"E3",X"DB",
		X"8B",X"E3",X"EF",X"8B",X"E3",X"2C",X"FB",X"DE",X"5C",X"63",X"FB",X"B7",X"00",X"97",X"57",X"FB",
		X"8F",X"B9",X"9D",X"FB",X"9A",X"5D",X"4D",X"5C",X"63",X"FB",X"0D",X"FB",X"9B",X"B2",X"C1",X"55",
		X"4D",X"97",X"BF",X"FF",X"96",X"E3",X"DB",X"0D",X"15",X"93",X"8B",X"B7",X"25",X"9F",X"D6",X"BF",
		X"9E",X"4D",X"5C",X"63",X"FB",X"0D",X"1D",X"B7",X"74",X"53",X"A3",X"C2",X"FC",X"A3",X"2A",X"FC",
		X"0D",X"15",X"1D",X"05",X"1C",X"61",X"41",X"40",X"EF",X"EF",X"EF",X"EF",X"8F",X"20",X"EF",X"98",
		X"20",X"EF",X"98",X"20",X"EF",X"DD",X"20",X"EF",X"DD",X"20",X"8B",X"DD",X"04",X"AB",X"EF",X"24",
		X"BF",X"EE",X"44",X"BF",X"00",X"64",X"8F",X"7B",X"F8",X"E0",X"68",X"FF",X"C1",X"8B",X"8B",X"E0",
		X"79",X"FF",X"C1",X"5C",X"8F",X"9B",X"5C",X"8F",X"9B",X"1C",X"97",X"75",X"FB",X"8F",X"EF",X"BD",
		X"5C",X"99",X"FF",X"1C",X"8A",X"40",X"29",X"09",X"1D",X"24",X"15",X"30",X"09",X"34",X"30",X"09",
		X"11",X"77",X"10",X"09",X"34",X"05",X"77",X"66",X"7E",X"5E",X"56",X"77",X"35",X"8A",X"8A",X"4C",
		X"D0",X"69",X"9B",X"E6",X"A3",X"9E",X"FC",X"1C",X"97",X"9A",X"DB",X"8F",X"A9",X"B9",X"5C",X"9C",
		X"FF",X"97",X"9D",X"D8",X"8F",X"99",X"B9",X"5C",X"5E",X"9B",X"1C",X"8A",X"58",X"65",X"45",X"45",
		X"45",X"45",X"45",X"45",X"41",X"8A",X"AA",X"61",X"75",X"75",X"75",X"75",X"75",X"75",X"69",X"8A",
		X"AA",X"6D",X"4D",X"4D",X"4D",X"4D",X"4D",X"4D",X"49",X"8A",X"5D",X"8A",X"8A",X"8F",X"C0",X"F8",
		X"C7",X"3D",X"A2",X"E0",X"F8",X"A3",X"C0",X"F8",X"A2",X"4A",X"FC",X"4B",X"3D",X"A2",X"B7",X"FC",
		X"4B",X"3D",X"FB",X"9F",X"5C",X"E0",X"DB",X"8F",X"9D",X"D8",X"E0",X"8B",X"63",X"AF",X"DF",X"E2",
		X"9F",X"A3",X"2F",X"F8",X"4D",X"97",X"9D",X"D8",X"8F",X"99",X"B9",X"5C",X"5E",X"9B",X"0D",X"8A",
		X"E0",X"4B",X"3D",X"E2",X"9A",X"5C",X"A6",X"BA",X"1C",X"53",X"8F",X"9D",X"D8",X"4C",X"C9",X"8B",
		X"4C",X"C9",X"8B",X"4C",X"C9",X"F8",X"8A",X"F9",X"8A",X"E0",X"5C",X"CA",X"DF",X"1C",X"97",X"B9",
		X"D8",X"B2",X"37",X"CB",X"B3",X"92",X"B2",X"70",X"BF",X"CB",X"B3",X"60",X"9B",X"34",X"53",X"B3",
		X"93",X"B3",X"1C",X"05",X"1A",X"41",X"8B",X"8A",X"E6",X"F3",X"DD",X"B5",X"F3",X"FD",X"B5",X"F0",
		X"D0",X"05",X"80",X"E1",X"FD",X"D4",X"15",X"F5",X"23",X"CC",X"F3",X"3D",X"B5",X"FF",X"37",X"15",
		X"D4",X"A6",X"2B",X"C2",X"8B",X"1E",X"45",X"5D",X"4D",X"01",X"10",X"73",X"57",X"89",X"2D",X"98",
		X"F6",X"2A",X"E0",X"46",X"51",X"53",X"53",X"B7",X"51",X"98",X"D2",X"98",X"D2",X"00",X"53",X"C1",
		X"8B",X"B7",X"64",X"8F",X"58",X"FC",X"97",X"B5",X"B5",X"9F",X"B7",X"BF",X"4C",X"27",X"8F",X"58",
		X"FC",X"97",X"BD",X"B5",X"9F",X"B7",X"BF",X"4C",X"27",X"E2",X"FF",X"A3",X"B8",X"B5",X"E2",X"DF",
		X"A3",X"DD",X"B5",X"A3",X"D8",X"B5",X"8F",X"43",X"FC",X"FB",X"FE",X"53",X"C1",X"8B",X"B7",X"64",
		X"A3",X"9F",X"B5",X"E6",X"A3",X"9F",X"B5",X"0D",X"1D",X"05",X"1C",X"98",X"45",X"98",X"03",X"0D",
		X"00",X"19",X"B7",X"C3",X"FB",X"9B",X"97",X"64",X"40",X"8F",X"42",X"FC",X"E0",X"4B",X"7D",X"CF",
		X"BE",X"96",X"B7",X"24",X"1C",X"10",X"ED",X"85",X"84",X"87",X"3E",X"4E",X"72",X"71",X"0D",X"53",
		X"53",X"87",X"98",X"1B",X"F0",X"8B",X"F1",X"10",X"88",X"F0",X"05",X"80",X"10",X"AF",X"80",X"69",
		X"2D",X"DB",X"DB",X"DB",X"8F",X"D8",X"BE",X"D0",X"DB",X"1B",X"F3",X"BF",X"D0",X"96",X"0C",X"19",
		X"88",X"BE",X"19",X"5E",X"BE",X"19",X"27",X"BE",X"19",X"0D",X"BE",X"19",X"93",X"9E",X"19",X"AC",
		X"BE",X"19",X"8C",X"BE",X"19",X"1E",X"9E",X"0D",X"15",X"1D",X"1C",X"0D",X"5C",X"97",X"9A",X"69",
		X"D2",X"8B",X"45",X"5C",X"97",X"9A",X"D9",X"05",X"8B",X"4D",X"5C",X"55",X"9E",X"DB",X"F3",X"BF",
		X"D0",X"8F",X"58",X"FC",X"96",X"A5",X"8B",X"E3",X"BF",X"15",X"19",X"C3",X"BE",X"0D",X"5C",X"97",
		X"9A",X"69",X"D2",X"8B",X"45",X"5C",X"97",X"9A",X"D8",X"8B",X"5C",X"97",X"9A",X"D9",X"05",X"8B",
		X"4D",X"DB",X"F3",X"BF",X"D0",X"8F",X"19",X"FC",X"96",X"85",X"8B",X"A5",X"15",X"19",X"C3",X"BE",
		X"0D",X"5C",X"97",X"9A",X"69",X"D2",X"8B",X"45",X"5C",X"97",X"9A",X"D8",X"8B",X"5C",X"97",X"9A",
		X"D9",X"05",X"8B",X"4D",X"45",X"DB",X"F3",X"BF",X"D0",X"8F",X"58",X"FC",X"96",X"4D",X"E0",X"8B",
		X"E8",X"C9",X"9E",X"FD",X"DC",X"0D",X"A5",X"8B",X"85",X"05",X"5C",X"55",X"9E",X"15",X"19",X"C3",
		X"BE",X"0D",X"5C",X"97",X"9A",X"69",X"D2",X"8B",X"45",X"5C",X"97",X"9A",X"D9",X"05",X"8B",X"4D",
		X"DB",X"F3",X"BF",X"D0",X"8F",X"58",X"FC",X"96",X"E0",X"26",X"AE",X"97",X"0D",X"5C",X"97",X"9A",
		X"D0",X"8B",X"5C",X"97",X"9A",X"D1",X"0D",X"81",X"8B",X"A1",X"19",X"C9",X"BE",X"15",X"93",X"93",
		X"19",X"C3",X"BE",X"0D",X"5C",X"97",X"9A",X"69",X"D2",X"8B",X"45",X"5C",X"97",X"9A",X"D9",X"8B",
		X"5C",X"97",X"9A",X"D8",X"05",X"8B",X"4D",X"45",X"DB",X"F3",X"BF",X"D0",X"8F",X"58",X"FC",X"96",
		X"53",X"62",X"AE",X"FB",X"C7",X"05",X"15",X"19",X"C3",X"BE",X"A4",X"69",X"2D",X"DB",X"DB",X"DB",
		X"DB",X"F3",X"BF",X"D0",X"8F",X"19",X"FC",X"96",X"F0",X"8B",X"F1",X"05",X"4D",X"DB",X"55",X"F3",
		X"BF",X"D0",X"8F",X"58",X"FC",X"96",X"15",X"B2",X"C1",X"93",X"A4",X"69",X"D2",X"A3",X"9F",X"DC",
		X"84",X"DB",X"55",X"F3",X"BF",X"D0",X"8F",X"58",X"FC",X"96",X"15",X"B2",X"93",X"D9",X"84",X"5C",
		X"55",X"9E",X"FE",X"A5",X"8B",X"E3",X"BF",X"8B",X"A2",X"9F",X"DC",X"C6",X"A3",X"9F",X"DC",X"AF",
		X"28",X"0D",X"A1",X"8A",X"81",X"15",X"19",X"C3",X"BE",X"0D",X"0D",X"A2",X"BB",X"DC",X"DB",X"DB",
		X"F3",X"BF",X"D0",X"8F",X"43",X"FC",X"96",X"F9",X"8B",X"F8",X"84",X"DB",X"F3",X"BF",X"D0",X"A2",
		X"BB",X"DC",X"45",X"E6",X"D9",X"DB",X"3F",X"45",X"FB",X"BF",X"5C",X"55",X"9E",X"8F",X"58",X"FC",
		X"05",X"DB",X"D0",X"F3",X"BF",X"96",X"A1",X"8B",X"A1",X"05",X"DB",X"DB",X"D0",X"8F",X"43",X"FC",
		X"96",X"E3",X"BF",X"19",X"C9",X"BE",X"97",X"BF",X"BF",X"4C",X"91",X"03",X"FC",X"97",X"9B",X"DF",
		X"4C",X"91",X"47",X"FC",X"1C",X"60",X"DE",X"35",X"45",X"5D",X"4D",X"55",X"97",X"F2",X"BA",X"DB",
		X"1B",X"D0",X"A0",X"78",X"BF",X"D1",X"B2",X"C9",X"93",X"B2",X"C8",X"53",X"15",X"0C",X"71",X"DF",
		X"71",X"DF",X"C6",X"B6",X"DB",X"79",X"DF",X"79",X"DF",X"E6",X"79",X"FF",X"EB",X"B5",X"79",X"B5",
		X"C8",X"A5",X"B6",X"F3",X"79",X"BB",X"79",X"9B",X"79",X"BB",X"79",X"FF",X"79",X"BB",X"EB",X"B5",
		X"79",X"B5",X"C8",X"A4",X"5C",X"09",X"9F",X"85",X"8B",X"A5",X"0D",X"1D",X"05",X"1C",X"BA",X"FA",
		X"BA",X"FE",X"9E",X"20",X"9E",X"04",X"BA",X"BA",X"BA",X"BE",X"9E",X"41",X"BA",X"FB",X"BA",X"FF",
		X"9E",X"45",X"9E",X"68",X"9E",X"25",X"9E",X"21",X"45",X"5D",X"55",X"4D",X"45",X"A2",X"B7",X"FC",
		X"60",X"9F",X"AF",X"BA",X"A2",X"97",X"FC",X"60",X"9F",X"AE",X"9B",X"05",X"B6",X"99",X"05",X"A3",
		X"9B",X"DC",X"D8",X"DB",X"DB",X"F3",X"BF",X"D0",X"8F",X"0E",X"BA",X"96",X"4D",X"8B",X"8B",X"F9",
		X"8B",X"E0",X"5D",X"4D",X"DB",X"DB",X"F3",X"BF",X"D0",X"8F",X"43",X"FC",X"96",X"E0",X"26",X"A6",
		X"DB",X"AF",X"9E",X"8B",X"E0",X"06",X"AE",X"FF",X"E2",X"9F",X"B6",X"9F",X"53",X"0D",X"1D",X"4B",
		X"0D",X"AE",X"FA",X"F0",X"8B",X"F1",X"8B",X"8B",X"E0",X"5C",X"73",X"BA",X"E2",X"9F",X"A3",X"9F",
		X"B5",X"0D",X"15",X"1D",X"05",X"1C",X"55",X"DB",X"DB",X"F3",X"BF",X"D0",X"8F",X"43",X"FC",X"96",
		X"A5",X"8B",X"85",X"8B",X"15",X"81",X"8B",X"A1",X"1C",X"B2",X"9A",X"9F",X"BF",X"90",X"9A",X"BB",
		X"BB",X"31",X"9A",X"BB",X"9F",X"9C",X"FE",X"BB",X"BF",X"C6",X"DE",X"BB",X"BF",X"DB",X"FA",X"BB",
		X"BF",X"83",X"FA",X"BB",X"BF",X"E0",X"FA",X"BB",X"BF",X"59",X"FA",X"BB",X"BF",X"BE",X"DA",X"BB",
		X"BF",X"98",X"DA",X"BB",X"BF",X"E9",X"DA",X"FB",X"BF",X"A0",X"DA",X"FF",X"BF",X"03",X"DA",X"9B",
		X"BF",X"71",X"DA",X"9B",X"BF",X"BF",X"B7",X"BB",X"BF",X"D7",X"B7",X"9F",X"BF",X"CB",X"B7",X"9B",
		X"9F",X"CD",X"B7",X"BB",X"9F",X"2E",X"B7",X"9F",X"9F",X"31",X"B7",X"BB",X"BB",X"41",X"B7",X"BB",
		X"BB",X"92",X"97",X"9F",X"BB",X"98",X"DA",X"9B",X"BF",X"9D",X"97",X"DF",X"BF",X"A0",X"DA",X"FF",
		X"BF",X"55",X"10",X"88",X"A0",X"10",X"AF",X"80",X"15",X"1C",X"D9",X"F8",X"DD",X"F9",X"F9",X"FD",
		X"F8",X"CD",X"F5",X"ED",X"FD",X"F8",X"BD",X"FD",X"CD",X"9D",X"FD",X"D9",X"BF",X"B0",X"EB",X"D8",
		X"B5",X"FD",X"02",X"B7",X"FD",X"EF",X"D8",X"E9",X"F8",X"DD",X"F9",X"CD",X"F9",X"FD",X"F8",X"ED",
		X"EC",X"BD",X"FD",X"CD",X"9D",X"FD",X"F9",X"AD",X"FD",X"CD",X"8D",X"FD",X"F9",X"BF",X"B0",X"9D",
		X"D8",X"B5",X"FD",X"DD",X"B7",X"ED",X"C6",X"D8",X"E9",X"FD",X"3F",X"DC",X"C8",X"EC",X"FD",X"FB",
		X"87",X"D8",X"F4",X"C0",X"C5",X"FD",X"45",X"B9",X"C9",X"87",X"FD",X"AB",X"D8",X"B4",X"FD",X"02",
		X"B6",X"FD",X"AB",X"D8",X"3F",X"9B",X"FC",X"BF",X"9F",X"BF",X"BF",X"9B",X"FD",X"BF",X"9F",X"BF",
		X"BF",X"AE",X"FC",X"BF",X"BB",X"BF",X"BF",X"9B",X"FD",X"BF",X"9F",X"BF",X"BF",X"9B",X"E6",X"BF",
		X"9F",X"BF",X"BF",X"9B",X"86",X"BF",X"9F",X"BF",X"BF",X"9B",X"A3",X"BF",X"9F",X"BF",X"BF",X"96",
		X"A7",X"BF",X"BB",X"BF",X"BF",X"96",X"A3",X"BF",X"96",X"BF",X"BF",X"9B",X"FC",X"BF",X"9F",X"BF",
		X"BF",X"9B",X"FD",X"BF",X"9F",X"BF",X"BF",X"96",X"FC",X"BF",X"FF",X"BF",X"BF",X"BA",X"86",X"BF",
		X"BB",X"BF",X"BF",X"BA",X"E6",X"BF",X"BB",X"BF",X"BF",X"BA",X"A7",X"BF",X"BB",X"BF",X"BF",X"AE",
		X"A3",X"BF",X"E9",X"C8",X"DF",X"2E",X"D8",X"C1",X"C0",X"E5",X"FD",X"D8",X"FD",X"65",X"FB",X"ED",
		X"A7",X"FD",X"04",X"D8",X"81",X"FD",X"02",X"83",X"FD",X"04",X"D8",X"3F",X"9B",X"36",X"BF",X"9F",
		X"BF",X"BF",X"9B",X"3E",X"BF",X"9F",X"BF",X"BF",X"AE",X"36",X"BF",X"BB",X"BF",X"BF",X"9B",X"3E",
		X"BF",X"9F",X"BF",X"BF",X"9B",X"A4",X"BF",X"9F",X"BF",X"BF",X"9B",X"A1",X"BF",X"9F",X"BF",X"BF",
		X"9B",X"CD",X"BF",X"9F",X"BF",X"BF",X"96",X"AD",X"BF",X"BB",X"BF",X"BF",X"96",X"CD",X"BF",X"96",
		X"BF",X"BF",X"9B",X"36",X"BF",X"9F",X"BF",X"BF",X"9B",X"3E",X"BF",X"9F",X"BF",X"BF",X"96",X"36",
		X"BF",X"FF",X"BF",X"BF",X"BA",X"A1",X"BF",X"BB",X"BF",X"BF",X"BA",X"A4",X"BF",X"BB",X"BF",X"BF",
		X"BA",X"AD",X"BF",X"BB",X"BF",X"BF",X"AE",X"CD",X"BF",X"D9",X"E8",X"FF",X"8F",X"EC",X"E1",X"BC",
		X"D1",X"FD",X"F9",X"FD",X"F8",X"FD",X"51",X"F9",X"FD",X"93",X"FD",X"A1",X"EC",X"A1",X"FD",X"02",
		X"A3",X"FD",X"A1",X"EC",X"3F",X"9B",X"B9",X"9F",X"9B",X"F1",X"9F",X"9B",X"A8",X"9F",X"9B",X"3F",
		X"9F",X"9B",X"73",X"9F",X"9B",X"6A",X"9F",X"9B",X"3C",X"9F",X"9B",X"2D",X"9F",X"9B",X"BF",X"BB",
		X"9B",X"AF",X"BB",X"9B",X"E6",X"BB",X"9B",X"AD",X"BB",X"9B",X"7F",X"BB",X"9B",X"6E",X"BB",X"9B",
		X"75",X"BB",X"9B",X"BF",X"9B",X"9B",X"EE",X"9B",X"9B",X"F4",X"9B",X"9B",X"75",X"BB",X"9B",X"BF",
		X"9B",X"9B",X"EE",X"9B",X"9B",X"6E",X"BB",X"9B",X"75",X"BB",X"9B",X"BF",X"9B",X"9B",X"7F",X"BB",
		X"9B",X"6E",X"BB",X"9B",X"75",X"BB",X"9B",X"AD",X"BB",X"9B",X"7F",X"BB",X"9B",X"6E",X"BB",X"9B",
		X"75",X"BB",X"9B",X"BF",X"9B",X"9B",X"EE",X"9B",X"9B",X"F4",X"9B",X"9B",X"37",X"9B",X"9B",X"3D",
		X"9B",X"9B",X"BF",X"FF",X"9B",X"BD",X"FF",X"9B",X"A4",X"FF",X"9B",X"3D",X"FF",X"9B",X"BE",X"DF",
		X"9B",X"B4",X"DF",X"9B",X"2E",X"DF",X"9B",X"BF",X"FB",X"9B",X"B4",X"FB",X"9B",X"B4",X"DF",X"9B",
		X"2E",X"DF",X"9B",X"BF",X"FB",X"9B",X"BE",X"DF",X"9B",X"B4",X"DF",X"9B",X"2E",X"DF",X"9B",X"3D",
		X"FF",X"9B",X"BE",X"DF",X"9B",X"B4",X"DF",X"9B",X"A4",X"FF",X"9B",X"3D",X"FF",X"9B",X"BE",X"DF",
		X"9B",X"B4",X"DF",X"9B",X"2E",X"DF",X"9B",X"BF",X"FB",X"9B",X"B4",X"FB",X"9B",X"26",X"FB",X"9B",
		X"AF",X"DB",X"9B",X"3F",X"DB",X"9B",X"BF",X"BE",X"9B",X"3F",X"BE",X"9B",X"25",X"BE",X"9B",X"3F",
		X"9E",X"9B",X"B7",X"BA",X"9B",X"27",X"BA",X"9B",X"B5",X"9A",X"9B",X"BF",X"FE",X"D9",X"C8",X"F9",
		X"FD",X"F8",X"CD",X"FF",X"94",X"CC",X"E1",X"F2",X"D1",X"FD",X"51",X"F9",X"FD",X"93",X"FD",X"B8",
		X"CC",X"A1",X"FD",X"02",X"A3",X"FD",X"B8",X"CC",X"3F",X"9F",X"73",X"9B",X"FF",X"BF",X"BF",X"9F",
		X"3C",X"9B",X"FF",X"BF",X"BF",X"9F",X"ED",X"9B",X"FF",X"BF",X"BF",X"9F",X"73",X"BB",X"FF",X"BF",
		X"BF",X"9F",X"3C",X"BB",X"FF",X"BF",X"BF",X"9F",X"ED",X"BB",X"FF",X"BF",X"BF",X"9F",X"73",X"9F",
		X"FF",X"BF",X"BF",X"9F",X"3C",X"9F",X"FF",X"BF",X"BF",X"9F",X"ED",X"9F",X"FF",X"BF",X"BF",X"9F",
		X"73",X"BF",X"FF",X"BF",X"BF",X"9F",X"3C",X"BF",X"FF",X"BF",X"BF",X"9F",X"ED",X"BF",X"FF",X"BF",
		X"BF",X"9F",X"A4",X"9F",X"9B",X"BF",X"BF",X"9F",X"2F",X"9F",X"9B",X"BF",X"BF",X"9F",X"98",X"9F",
		X"9B",X"BF",X"BF",X"9F",X"A4",X"BF",X"9B",X"BF",X"BF",X"9F",X"2F",X"BF",X"9B",X"BF",X"BF",X"9F",
		X"98",X"BF",X"9F",X"B0",X"9F",X"BB",X"BF",X"BF",X"9F",X"A4",X"9F",X"BB",X"BF",X"BF",X"9F",X"A3",
		X"9F",X"BB",X"BF",X"BF",X"9F",X"B0",X"BF",X"BB",X"BF",X"BF",X"9F",X"A4",X"BF",X"BB",X"BF",X"BF",
		X"9F",X"A3",X"BF",X"BB",X"BF",X"BF",X"9F",X"E6",X"9F",X"9F",X"BF",X"BF",X"9F",X"B5",X"9F",X"9F",
		X"BF",X"BF",X"9F",X"F2",X"9F",X"9F",X"BF",X"BF",X"9F",X"E6",X"BF",X"9F",X"BF",X"BF",X"9F",X"B5",
		X"BF",X"9F",X"BF",X"BF",X"9F",X"F2",X"BF",X"D9",X"EC",X"E9",X"EC",X"F8",X"CD",X"D8",X"ED",X"DD",
		X"FD",X"F9",X"FD",X"CD",X"FD",X"FD",X"F7",X"ED",X"F7",X"F5",X"D5",X"B5",X"FD",X"02",X"BD",X"FD",
		X"ED",X"AD",X"FD",X"D9",X"B7",X"FD",X"D0",X"E8",X"99",X"FD",X"02",X"A9",X"FD",X"02",X"AB",X"FD",
		X"C5",X"E8",X"3F",X"D9",X"C8",X"E9",X"C8",X"DC",X"C8",X"D1",X"D9",X"F9",X"FD",X"F8",X"C9",X"D8",
		X"C9",X"EC",X"CD",X"FD",X"F7",X"DD",X"FD",X"ED",X"D7",X"CD",X"FD",X"C9",X"F3",X"FC",X"FD",X"F5",
		X"D5",X"B5",X"FD",X"02",X"BD",X"7D",X"02",X"AD",X"7D",X"02",X"89",X"7D",X"02",X"B7",X"FD",X"95",
		X"E8",X"91",X"FD",X"02",X"93",X"FD",X"99",X"E8",X"FD",X"7D",X"DD",X"D9",X"B5",X"FD",X"DD",X"AD",
		X"FD",X"F8",X"89",X"FD",X"F8",X"B7",X"CD",X"AE",X"E8",X"E9",X"FD",X"DC",X"FD",X"3F",X"D9",X"EC",
		X"DD",X"DD",X"F9",X"FD",X"F8",X"E9",X"E9",X"EC",X"CD",X"DD",X"D8",X"CD",X"DC",X"EC",X"FC",X"DD",
		X"EC",X"ED",X"F5",X"E0",X"D1",X"CD",X"FD",X"FF",X"B5",X"FD",X"2E",X"ED",X"DF",X"C9",X"FB",X"BD",
		X"FD",X"E9",X"AD",X"FD",X"E9",X"89",X"FD",X"E9",X"B5",X"FD",X"DD",X"B7",X"E0",X"40",X"E8",X"99",
		X"7D",X"22",X"A9",X"7D",X"22",X"9C",X"7D",X"22",X"B5",X"FD",X"CD",X"91",X"FD",X"02",X"93",X"FD",
		X"74",X"E8",X"E9",X"FD",X"DC",X"FD",X"3F",X"D9",X"C9",X"FD",X"FD",X"DD",X"FC",X"F9",X"FD",X"F8",
		X"CD",X"ED",X"ED",X"CD",X"FD",X"E9",X"C9",X"D8",X"CD",X"C9",X"C8",X"FC",X"FD",X"DC",X"C9",X"EC",
		X"CD",X"F5",X"82",X"BD",X"FD",X"FC",X"AD",X"FD",X"ED",X"89",X"FD",X"06",X"B5",X"FD",X"02",X"B7",
		X"FD",X"1B",X"E8",X"9D",X"FD",X"26",X"8D",X"FD",X"36",X"BC",X"FD",X"ED",X"B5",X"FD",X"DD",X"B7",
		X"82",X"13",X"E8",X"E9",X"FD",X"DC",X"FD",X"3F",X"D9",X"F8",X"FD",X"7F",X"DD",X"FD",X"F9",X"FD",
		X"F8",X"CD",X"E9",X"F8",X"ED",X"7A",X"CD",X"FD",X"D8",X"CD",X"DC",X"F8",X"C9",X"67",X"FC",X"FD",
		X"EC",X"CD",X"D1",X"DB",X"F5",X"F8",X"B5",X"FD",X"02",X"BD",X"FD",X"06",X"AD",X"FD",X"06",X"89",
		X"FD",X"06",X"B7",X"FD",X"EB",X"C8",X"BD",X"FD",X"E5",X"AD",X"FD",X"E5",X"89",X"FD",X"E5",X"91",
		X"FD",X"02",X"93",X"FD",X"EF",X"C8",X"E9",X"FD",X"DC",X"FD",X"3F",X"D9",X"E8",X"FD",X"FD",X"DD",
		X"DD",X"F9",X"FD",X"F8",X"FD",X"BD",X"FD",X"F7",X"BF",X"37",X"85",X"C8",X"FD",X"FD",X"9D",X"FD",
		X"D9",X"9F",X"C9",X"85",X"C8",X"3F",X"D9",X"CD",X"FD",X"C9",X"DD",X"C9",X"F9",X"DD",X"F8",X"FD",
		X"F5",X"CD",X"B5",X"FD",X"02",X"B7",X"FD",X"B3",X"C8",X"3F",X"FD",X"FF",X"DD",X"DD",X"F9",X"DD",
		X"F8",X"CD",X"D9",X"F8",X"F5",X"CC",X"BD",X"FD",X"F5",X"B5",X"FD",X"02",X"B7",X"FD",X"69",X"C8",
		X"9D",X"FD",X"DD",X"F5",X"D9",X"9F",X"D9",X"69",X"C8",X"F5",X"E4",X"DD",X"DD",X"FD",X"3F",X"BD",
		X"FD",X"36",X"B5",X"FD",X"02",X"B7",X"FD",X"40",X"C8",X"9D",X"FD",X"02",X"F5",X"02",X"9F",X"FD",
		X"40",X"C8",X"3F",X"D9",X"E8",X"F8",X"ED",X"D1",X"F9",X"F9",X"FD",X"DD",X"DD",X"FD",X"CF",X"F5",
		X"E5",X"B5",X"FD",X"02",X"BD",X"FD",X"37",X"99",X"7D",X"02",X"B7",X"FD",X"1D",X"C8",X"91",X"FD",
		X"02",X"93",X"FD",X"46",X"C8",X"3F",X"D9",X"C8",X"F8",X"CD",X"D1",X"F9",X"F5",X"E9",X"FD",X"3D",
		X"DD",X"DD",X"F9",X"FD",X"B5",X"FD",X"02",X"B7",X"FD",X"2F",X"C8",X"B5",X"FD",X"DD",X"99",X"FD",
		X"02",X"BD",X"FD",X"E9",X"B7",X"E9",X"1A",X"C8",X"91",X"FD",X"02",X"93",X"FD",X"24",X"C8",X"3F",
		X"FD",X"BF",X"DD",X"ED",X"F9",X"FD",X"D9",X"D8",X"F8",X"F9",X"BD",X"FD",X"ED",X"99",X"7D",X"02",
		X"BF",X"77",X"F8",X"F5",X"3F",X"FD",X"80",X"DD",X"FD",X"F9",X"FD",X"D9",X"C8",X"F8",X"FD",X"B8",
		X"FD",X"DD",X"BA",X"C8",X"C0",X"F5",X"3F",X"E9",X"F8",X"D8",X"FD",X"DF",X"9D",X"F5",X"C1",X"EC",
		X"E5",X"FD",X"65",X"FB",X"ED",X"A7",X"FD",X"F3",X"F5",X"81",X"FD",X"02",X"83",X"FD",X"F3",X"F5",
		X"3F",X"BB",X"A4",X"BF",X"9F",X"BF",X"BF",X"BB",X"36",X"BF",X"9F",X"BF",X"BF",X"BB",X"47",X"BF",
		X"9F",X"BF",X"BF",X"FB",X"2D",X"9F",X"FB",X"BF",X"BF",X"FF",X"73",X"9F",X"BB",X"BF",X"BF",X"BA",
		X"2D",X"9F",X"B3",X"BF",X"BF",X"CD",X"DD",X"D8",X"FD",X"E9",X"DD",X"ED",X"7D",X"D5",X"F8",X"95",
		X"FD",X"02",X"AD",X"FD",X"03",X"A9",X"7D",X"FD",X"98",X"FD",X"DD",X"97",X"FD",X"8A",X"F5",X"E9",
		X"DD",X"ED",X"7F",X"95",X"FD",X"DD",X"AD",X"FD",X"03",X"A9",X"7D",X"FD",X"98",X"FD",X"DD",X"97",
		X"F8",X"59",X"F5",X"E9",X"DD",X"ED",X"3D",X"95",X"FD",X"02",X"AD",X"FD",X"03",X"A9",X"7D",X"FD",
		X"98",X"FD",X"DD",X"97",X"FD",X"41",X"F5",X"3F",X"E9",X"CD",X"ED",X"D9",X"CD",X"CD",X"D8",X"CD",
		X"D5",X"C9",X"95",X"FD",X"02",X"A9",X"7D",X"FD",X"AD",X"7D",X"ED",X"8D",X"7D",X"02",X"97",X"FD",
		X"73",X"F5",X"D8",X"ED",X"95",X"FD",X"DD",X"A9",X"7D",X"02",X"AD",X"FD",X"7A",X"97",X"FC",X"2D",
		X"F5",X"3F",X"DC",X"EC",X"EC",X"F9",X"C9",X"3D",X"FC",X"FD",X"F1",X"F3",X"B1",X"FD",X"02",X"89",
		X"FD",X"ED",X"BC",X"F5",X"FD",X"B3",X"FD",X"24",X"F5",X"B1",X"FD",X"DD",X"89",X"3D",X"02",X"BC",
		X"FD",X"02",X"B3",X"F3",X"1E",X"F5",X"3F",X"FC",X"FD",X"EC",X"CD",X"F1",X"CD",X"C9",X"E0",X"C5",
		X"F8",X"DC",X"C8",X"89",X"FD",X"32",X"9C",X"FD",X"02",X"85",X"FD",X"02",X"87",X"FD",X"D9",X"D5",
		X"B1",X"FD",X"02",X"89",X"FD",X"BF",X"B3",X"FD",X"02",X"F5",X"3F",X"C9",X"7D",X"FC",X"DD",X"DC",
		X"CD",X"EC",X"FD",X"F1",X"CD",X"89",X"BD",X"FD",X"B1",X"FD",X"02",X"B3",X"FD",X"CF",X"D5",X"FC",
		X"FC",X"C9",X"7D",X"89",X"FD",X"F9",X"BC",X"3D",X"02",X"B1",X"FD",X"DD",X"B3",X"F4",X"D3",X"D5",
		X"3F",X"D9",X"FD",X"3F",X"4D",X"8F",X"91",X"97",X"97",X"1A",X"9E",X"9F",X"F3",X"D3",X"10",X"ED",
		X"91",X"59",X"65",X"10",X"F7",X"C0",X"72",X"4A",X"2D",X"72",X"FB",X"2D",X"6E",X"72",X"CB",X"2D",
		X"72",X"75",X"34",X"72",X"65",X"0D",X"98",X"44",X"5C",X"61",X"9F",X"5C",X"63",X"DB",X"00",X"FB",
		X"9F",X"5D",X"97",X"0E",X"97",X"5C",X"F0",X"96",X"97",X"CF",X"A2",X"8F",X"3A",X"99",X"5C",X"9C",
		X"FF",X"97",X"26",X"97",X"8F",X"98",X"B9",X"5C",X"9C",X"FF",X"97",X"14",X"97",X"8F",X"25",X"B9",
		X"5C",X"9C",X"FF",X"FB",X"BE",X"8F",X"41",X"F9",X"E3",X"BF",X"8A",X"B7",X"00",X"8B",X"1D",X"B4",
		X"D6",X"F3",X"BF",X"96",X"F5",X"D4",X"19",X"E0",X"B3",X"8A",X"79",X"25",X"1D",X"15",X"01",X"29",
		X"09",X"10",X"24",X"1D",X"11",X"10",X"8A",X"8A",X"25",X"05",X"10",X"1D",X"30",X"05",X"25",X"77",
		X"24",X"05",X"10",X"24",X"6B",X"8A",X"AA",X"24",X"09",X"77",X"05",X"3C",X"05",X"11",X"04",X"24",
		X"05",X"77",X"24",X"05",X"10",X"24",X"6B",X"8A",X"8A",X"8A",X"51",X"6A",X"77",X"56",X"77",X"77",
		X"11",X"04",X"30",X"30",X"05",X"29",X"24",X"77",X"10",X"05",X"24",X"24",X"1D",X"29",X"01",X"10",
		X"8A",X"AA",X"6A",X"77",X"72",X"77",X"77",X"10",X"24",X"15",X"24",X"1D",X"11",X"77",X"30",X"15",
		X"0D",X"8A",X"AA",X"6A",X"77",X"52",X"77",X"77",X"05",X"34",X"30",X"09",X"0D",X"10",X"8A",X"AA",
		X"6A",X"77",X"66",X"77",X"77",X"11",X"09",X"29",X"20",X"05",X"30",X"01",X"05",X"29",X"11",X"05",
		X"8A",X"AA",X"6A",X"77",X"46",X"77",X"77",X"2D",X"05",X"20",X"05",X"2D",X"10",X"8A",X"AA",X"6A",
		X"77",X"62",X"77",X"77",X"10",X"09",X"04",X"29",X"25",X"10",X"8A",X"AA",X"6A",X"77",X"42",X"77",
		X"77",X"31",X"04",X"24",X"24",X"09",X"29",X"10",X"8A",X"AA",X"6A",X"77",X"7E",X"77",X"77",X"05",
		X"3C",X"1D",X"24",X"8A",X"8A",X"DF",X"8A",X"A4",X"4B",X"AF",X"8B",X"FB",X"BE",X"8F",X"41",X"F9",
		X"B6",X"F6",X"A3",X"3D",X"B5",X"A2",X"BF",X"B5",X"D4",X"F5",X"18",X"D9",X"AE",X"49",X"18",X"D0",
		X"AF",X"D3",X"FF",X"8B",X"A4",X"60",X"9E",X"AF",X"DF",X"FB",X"9F",X"8F",X"25",X"F9",X"53",X"B3",
		X"E3",X"FF",X"5D",X"FB",X"A5",X"5C",X"64",X"BB",X"1D",X"A2",X"BD",X"B5",X"18",X"C1",X"AF",X"31",
		X"A4",X"60",X"9F",X"38",X"48",X"B3",X"60",X"BB",X"38",X"A2",X"F7",X"60",X"9B",X"38",X"DE",X"D7",
		X"60",X"FF",X"38",X"77",X"D7",X"60",X"DF",X"38",X"6A",X"D7",X"60",X"FB",X"38",X"D3",X"D3",X"60",
		X"DB",X"38",X"FF",X"B6",X"60",X"BE",X"AE",X"60",X"5C",X"62",X"B3",X"19",X"85",X"97",X"45",X"5D",
		X"97",X"71",X"B3",X"8F",X"DB",X"BD",X"5C",X"99",X"FF",X"A2",X"BD",X"B5",X"A3",X"3D",X"B5",X"18",
		X"C1",X"AF",X"61",X"1D",X"05",X"1C",X"8A",X"5D",X"24",X"1D",X"3C",X"05",X"77",X"09",X"24",X"8A",
		X"55",X"77",X"3D",X"11",X"29",X"04",X"34",X"8A",X"5D",X"77",X"24",X"1D",X"3D",X"8A",X"8A",X"5D",
		X"53",X"5C",X"FC",X"BB",X"E2",X"9E",X"5C",X"23",X"BB",X"5C",X"00",X"DF",X"97",X"4F",X"93",X"8F",
		X"6B",X"B9",X"5C",X"9C",X"FF",X"97",X"71",X"B3",X"8F",X"DB",X"BD",X"5C",X"99",X"FF",X"97",X"63",
		X"93",X"8F",X"37",X"99",X"5C",X"99",X"FF",X"97",X"3D",X"93",X"8F",X"A5",X"B9",X"5C",X"9C",X"FF",
		X"97",X"75",X"93",X"8F",X"23",X"B9",X"5C",X"9C",X"FF",X"97",X"20",X"93",X"8F",X"47",X"B9",X"5C",
		X"9C",X"FF",X"A2",X"BD",X"B5",X"69",X"3F",X"8F",X"7C",X"B9",X"97",X"B6",X"F7",X"AE",X"9B",X"97",
		X"8E",X"F7",X"5C",X"9C",X"FF",X"A3",X"3D",X"B5",X"A2",X"3F",X"B5",X"69",X"C2",X"D8",X"8F",X"B5",
		X"99",X"FB",X"FB",X"DA",X"97",X"FA",X"F7",X"A7",X"9B",X"97",X"93",X"F7",X"4D",X"5C",X"9C",X"FF",
		X"0D",X"8B",X"B7",X"48",X"84",X"69",X"9B",X"68",X"9B",X"79",X"83",X"A3",X"27",X"B9",X"84",X"69",
		X"F6",X"68",X"F6",X"DA",X"DA",X"D8",X"79",X"87",X"A3",X"33",X"BD",X"FE",X"9D",X"8F",X"83",X"B9",
		X"E3",X"90",X"8F",X"93",X"B9",X"97",X"2D",X"40",X"E2",X"D4",X"5C",X"C7",X"FF",X"E2",X"BE",X"17",
		X"AE",X"FB",X"D9",X"E2",X"F4",X"5C",X"C7",X"FF",X"E3",X"F0",X"A2",X"BD",X"B5",X"18",X"C1",X"AF",
		X"17",X"1D",X"19",X"85",X"97",X"8A",X"79",X"11",X"09",X"29",X"21",X"1D",X"01",X"04",X"30",X"15",
		X"24",X"1D",X"09",X"29",X"8A",X"8A",X"8A",X"61",X"56",X"72",X"52",X"66",X"46",X"62",X"8A",X"8A",
		X"8A",X"5D",X"2D",X"1D",X"20",X"05",X"10",X"77",X"34",X"05",X"30",X"77",X"11",X"30",X"05",X"25",
		X"1D",X"24",X"8A",X"8A",X"25",X"1D",X"21",X"21",X"1D",X"11",X"04",X"2D",X"24",X"1C",X"77",X"2D",
		X"05",X"20",X"05",X"2D",X"8A",X"AA",X"05",X"15",X"10",X"1C",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"3D",X"15",X"30",X"25",X"8A",X"8A",X"15",X"24",X"24",X"30",X"15",X"11",
		X"24",X"77",X"0D",X"09",X"25",X"05",X"77",X"10",X"09",X"04",X"29",X"25",X"8A",X"8A",X"09",X"29",
		X"77",X"8A",X"8A",X"09",X"21",X"21",X"8A",X"8A",X"8A",X"65",X"77",X"24",X"15",X"31",X"2D",X"05",
		X"77",X"0D",X"09",X"25",X"05",X"2D",X"77",X"8A",X"8A",X"8A",X"65",X"04",X"34",X"30",X"1D",X"01",
		X"3D",X"24",X"77",X"0D",X"09",X"25",X"05",X"2D",X"8A",X"8A",X"5D",X"97",X"4B",X"F7",X"5C",X"F0",
		X"96",X"8F",X"BF",X"BD",X"97",X"27",X"FC",X"5C",X"48",X"F7",X"8F",X"BF",X"FD",X"93",X"5C",X"48",
		X"F7",X"8F",X"BF",X"FC",X"93",X"5C",X"48",X"F7",X"9F",X"27",X"FC",X"E2",X"9B",X"8F",X"A5",X"99",
		X"97",X"43",X"F7",X"45",X"4D",X"5C",X"9C",X"FF",X"55",X"97",X"55",X"F7",X"BA",X"69",X"DA",X"AE",
		X"9B",X"97",X"29",X"F7",X"5C",X"9C",X"FF",X"97",X"BD",X"40",X"96",X"15",X"5C",X"9C",X"FF",X"55",
		X"97",X"55",X"F7",X"BA",X"69",X"25",X"AE",X"9B",X"97",X"29",X"F7",X"5C",X"9C",X"FF",X"15",X"0D",
		X"8B",X"8B",X"05",X"9B",X"C6",X"AF",X"7C",X"97",X"71",X"B3",X"8F",X"DB",X"BD",X"5C",X"99",X"FF",
		X"5C",X"62",X"B3",X"1D",X"19",X"85",X"97",X"8A",X"79",X"10",X"24",X"15",X"24",X"1D",X"11",X"77",
		X"30",X"15",X"0D",X"8A",X"5D",X"8A",X"8A",X"66",X"19",X"77",X"8A",X"8A",X"66",X"29",X"77",X"8A",
		X"8A",X"66",X"2D",X"77",X"8A",X"8A",X"66",X"34",X"77",X"8A",X"8A",X"66",X"0D",X"77",X"8A",X"8A",
		X"66",X"30",X"77",X"8A",X"8A",X"8A",X"65",X"09",X"19",X"77",X"77",X"77",X"77",X"77",X"8A",X"5D",
		X"8A",X"8A",X"8A",X"71",X"29",X"09",X"24",X"77",X"09",X"19",X"77",X"8A",X"5D",X"8A",X"8A",X"53",
		X"9F",X"FF",X"BF",X"4D",X"5D",X"45",X"F8",X"C1",X"6A",X"08",X"63",X"C1",X"08",X"85",X"05",X"8B",
		X"B7",X"01",X"1D",X"DE",X"AF",X"68",X"0D",X"C6",X"60",X"60",X"AF",X"6D",X"1C",X"5D",X"97",X"B5",
		X"D7",X"5C",X"F0",X"96",X"8F",X"BF",X"AF",X"9F",X"D2",X"60",X"5C",X"CC",X"D7",X"45",X"8F",X"BF",
		X"BF",X"9F",X"AF",X"BF",X"5C",X"CC",X"D7",X"9F",X"60",X"C2",X"97",X"8D",X"D7",X"8F",X"37",X"B9",
		X"5C",X"E1",X"D7",X"9F",X"40",X"C2",X"97",X"E9",X"D7",X"8F",X"13",X"B9",X"05",X"5C",X"E1",X"D7",
		X"97",X"71",X"B3",X"8F",X"DB",X"BD",X"5C",X"99",X"FF",X"5C",X"62",X"B3",X"1D",X"19",X"85",X"97",
		X"8A",X"79",X"05",X"34",X"30",X"09",X"0D",X"77",X"11",X"3D",X"05",X"11",X"19",X"8A",X"5D",X"8A",
		X"8A",X"04",X"72",X"77",X"8A",X"8A",X"8A",X"5D",X"04",X"52",X"77",X"8A",X"8A",X"53",X"7B",X"8B",
		X"B7",X"64",X"DE",X"AF",X"04",X"1C",X"45",X"5C",X"9C",X"FF",X"BA",X"1D",X"97",X"55",X"F7",X"26",
		X"AE",X"FF",X"97",X"29",X"F7",X"A4",X"45",X"5C",X"9C",X"FF",X"E2",X"9F",X"A3",X"BF",X"FC",X"05",
		X"5C",X"0C",X"9B",X"1C",X"5D",X"5C",X"00",X"DF",X"E2",X"9E",X"5C",X"23",X"BB",X"E2",X"D2",X"5C",
		X"4E",X"BB",X"FB",X"F2",X"5C",X"9E",X"9B",X"5C",X"62",X"B3",X"1D",X"19",X"85",X"97",X"5D",X"53",
		X"A3",X"FB",X"FC",X"97",X"6A",X"FC",X"8F",X"4E",X"FC",X"E6",X"B3",X"C1",X"55",X"4D",X"97",X"4F",
		X"F3",X"5C",X"F0",X"96",X"97",X"CF",X"A2",X"8F",X"3A",X"99",X"5C",X"9C",X"FF",X"97",X"67",X"F3",
		X"8F",X"98",X"B9",X"5C",X"9C",X"FF",X"97",X"75",X"F3",X"8F",X"55",X"B9",X"5C",X"9C",X"FF",X"97",
		X"60",X"F3",X"8F",X"DF",X"BD",X"5C",X"99",X"FF",X"0D",X"15",X"B2",X"4D",X"8F",X"57",X"9D",X"5C",
		X"4B",X"9B",X"0D",X"FB",X"A5",X"5C",X"64",X"BB",X"A3",X"3D",X"B5",X"A2",X"BD",X"B5",X"18",X"C1",
		X"AE",X"EE",X"A2",X"BF",X"B5",X"18",X"D9",X"AE",X"FB",X"18",X"D0",X"AE",X"B7",X"B6",X"0C",X"E7",
		X"B2",X"79",X"9F",X"CB",X"60",X"AF",X"AF",X"BB",X"53",X"C1",X"B3",X"B6",X"5C",X"C7",X"B2",X"71",
		X"9F",X"CB",X"60",X"16",X"AF",X"DF",X"E2",X"93",X"C1",X"E2",X"96",X"B3",X"B6",X"66",X"B2",X"A3",
		X"DB",X"DC",X"E0",X"A3",X"FB",X"DC",X"4B",X"38",X"0F",X"F3",X"60",X"9F",X"AE",X"B6",X"C6",X"D9",
		X"A2",X"3F",X"B5",X"69",X"F6",X"68",X"F6",X"DA",X"DA",X"E6",X"D8",X"E2",X"9F",X"1F",X"B7",X"44",
		X"60",X"B7",X"A6",X"BB",X"E2",X"DA",X"A3",X"BE",X"DC",X"53",X"A3",X"2F",X"F8",X"A3",X"76",X"FC",
		X"A3",X"B7",X"FC",X"E6",X"A3",X"FF",X"DC",X"A3",X"BD",X"FC",X"A3",X"82",X"FC",X"55",X"4D",X"5C",
		X"56",X"EF",X"5C",X"00",X"DF",X"97",X"71",X"B3",X"8F",X"DB",X"BD",X"5C",X"99",X"FF",X"97",X"0D",
		X"F3",X"8F",X"CF",X"BD",X"5C",X"99",X"FF",X"A3",X"3D",X"B5",X"A2",X"BD",X"B5",X"18",X"C1",X"AE",
		X"9A",X"A2",X"BF",X"B5",X"CA",X"69",X"DA",X"AE",X"68",X"5C",X"C0",X"8A",X"0D",X"15",X"19",X"66",
		X"D7",X"1D",X"19",X"85",X"97",X"8A",X"79",X"2D",X"05",X"20",X"05",X"2D",X"77",X"11",X"3D",X"05",
		X"11",X"19",X"8A",X"8A",X"2D",X"05",X"20",X"05",X"2D",X"77",X"29",X"04",X"0D",X"31",X"05",X"30",
		X"6B",X"8A",X"AA",X"24",X"09",X"77",X"10",X"05",X"24",X"04",X"34",X"77",X"2D",X"05",X"20",X"05",
		X"2D",X"6B",X"8A",X"8A",X"8A",X"51",X"2D",X"05",X"20",X"05",X"2D",X"77",X"29",X"09",X"7A",X"8A",
		X"8A",X"8A",X"5D",X"1C",X"15",X"2D",X"34",X"77",X"09",X"24",X"8A",X"65",X"77",X"19",X"11",X"1D",
		X"24",X"10",X"1C",X"09",X"39",X"8A",X"5D",X"77",X"05",X"20",X"09",X"0D",X"8A",X"8A",X"8A",X"59",
		X"24",X"1D",X"3C",X"05",X"77",X"09",X"24",X"77",X"76",X"77",X"2D",X"05",X"20",X"05",X"2D",X"77",
		X"34",X"04",X"24",X"05",X"10",X"8A",X"8A",X"5D",X"5C",X"63",X"DB",X"97",X"6A",X"FC",X"8F",X"4E",
		X"FC",X"53",X"A3",X"FB",X"FC",X"E6",X"B3",X"C1",X"55",X"4D",X"97",X"0A",X"D3",X"5C",X"F0",X"96",
		X"97",X"CF",X"A2",X"8F",X"3A",X"99",X"5C",X"9C",X"FF",X"97",X"22",X"D3",X"8F",X"98",X"B9",X"5C",
		X"9C",X"FF",X"97",X"74",X"D3",X"8F",X"55",X"B9",X"5C",X"9C",X"FF",X"97",X"0C",X"D3",X"8F",X"9B",
		X"BD",X"5C",X"99",X"FF",X"0D",X"15",X"B2",X"4D",X"8F",X"57",X"9D",X"5C",X"4B",X"9B",X"0D",X"FB",
		X"A5",X"5C",X"64",X"BB",X"A3",X"3D",X"B5",X"A2",X"BD",X"B5",X"18",X"C1",X"AE",X"EE",X"A2",X"BF",
		X"B5",X"18",X"D9",X"AE",X"FB",X"18",X"D0",X"AE",X"B7",X"B6",X"0C",X"E7",X"B2",X"79",X"9F",X"CB",
		X"60",X"EF",X"AF",X"BB",X"53",X"C1",X"B3",X"B6",X"5C",X"C7",X"B2",X"71",X"9F",X"CB",X"60",X"16",
		X"AF",X"DF",X"E2",X"D3",X"C1",X"E2",X"8B",X"B3",X"B6",X"66",X"E0",X"4B",X"AE",X"FB",X"C6",X"5C",
		X"A6",X"BA",X"B6",X"23",X"5C",X"63",X"DB",X"1D",X"19",X"85",X"97",X"8A",X"79",X"10",X"09",X"04",
		X"29",X"25",X"77",X"11",X"3D",X"05",X"11",X"19",X"8A",X"8A",X"10",X"09",X"04",X"29",X"25",X"77",
		X"29",X"04",X"0D",X"31",X"05",X"30",X"6B",X"8A",X"AA",X"24",X"09",X"77",X"05",X"3C",X"05",X"11",
		X"04",X"24",X"05",X"77",X"10",X"09",X"04",X"29",X"25",X"6B",X"8A",X"8A",X"8A",X"51",X"10",X"09",
		X"04",X"29",X"25",X"77",X"29",X"09",X"7A",X"8A",X"8A",X"8A",X"59",X"24",X"1D",X"3C",X"05",X"77",
		X"09",X"24",X"77",X"76",X"77",X"25",X"29",X"04",X"09",X"10",X"77",X"05",X"24",X"04",X"11",X"05",
		X"3C",X"05",X"8A",X"8A",X"5D",X"97",X"3A",X"B6",X"5C",X"F0",X"96",X"97",X"32",X"B6",X"8F",X"B8",
		X"99",X"5C",X"9C",X"FF",X"97",X"4D",X"B6",X"8F",X"B5",X"99",X"5C",X"9C",X"FF",X"97",X"FA",X"96",
		X"8F",X"B7",X"9D",X"5C",X"9C",X"FF",X"97",X"71",X"B3",X"8F",X"DB",X"BD",X"5C",X"99",X"FF",X"53",
		X"A3",X"B0",X"B5",X"FB",X"FF",X"97",X"7B",X"B6",X"8F",X"F1",X"B5",X"B2",X"C1",X"93",X"8B",X"B7",
		X"20",X"A2",X"BD",X"B5",X"D0",X"CA",X"69",X"DA",X"D8",X"A2",X"BF",X"B5",X"D1",X"CA",X"69",X"DA",
		X"D9",X"18",X"A8",X"AF",X"BB",X"18",X"2D",X"18",X"A0",X"AF",X"BB",X"18",X"0D",X"A4",X"07",X"E2",
		X"BA",X"AF",X"9F",X"53",X"A3",X"B0",X"B5",X"A3",X"3D",X"B5",X"A4",X"8F",X"B5",X"D9",X"5C",X"BD",
		X"96",X"84",X"8F",X"B7",X"DD",X"5C",X"BD",X"96",X"A2",X"BD",X"B5",X"18",X"C1",X"AF",X"39",X"5C",
		X"63",X"DB",X"1D",X"19",X"85",X"97",X"BB",X"9F",X"BF",X"BF",X"8A",X"79",X"31",X"04",X"24",X"24",
		X"09",X"29",X"77",X"11",X"3D",X"05",X"11",X"19",X"8A",X"8A",X"8A",X"5D",X"77",X"77",X"77",X"25",
		X"05",X"34",X"30",X"05",X"10",X"10",X"05",X"25",X"77",X"31",X"04",X"24",X"24",X"09",X"29",X"10",
		X"8A",X"AA",X"77",X"77",X"77",X"15",X"30",X"05",X"77",X"3D",X"1D",X"01",X"3D",X"2D",X"1D",X"01",
		X"3D",X"24",X"05",X"25",X"6B",X"8A",X"AA",X"8A",X"AA",X"8A",X"71",X"34",X"2D",X"15",X"1C",X"05",
		X"30",X"77",X"56",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"34",X"2D",X"15",X"1C",X"05",
		X"30",X"77",X"72",X"8A",X"8A",X"8A",X"69",X"04",X"34",X"8A",X"AA",X"8A",X"AA",X"2D",X"05",X"21",
		X"24",X"8A",X"AA",X"8A",X"AA",X"30",X"1D",X"01",X"3D",X"24",X"8A",X"AA",X"8A",X"AA",X"25",X"09",
		X"00",X"29",X"8A",X"AA",X"8A",X"AA",X"11",X"09",X"1D",X"29",X"1D",X"29",X"8A",X"8A",X"8A",X"69",
		X"77",X"77",X"77",X"77",X"04",X"34",X"8A",X"AA",X"8A",X"AA",X"77",X"77",X"2D",X"05",X"21",X"24",
		X"8A",X"AA",X"8A",X"AA",X"77",X"30",X"1D",X"01",X"3D",X"24",X"8A",X"AA",X"8A",X"AA",X"77",X"77",
		X"25",X"09",X"00",X"29",X"8A",X"AA",X"8A",X"AA",X"77",X"34",X"04",X"29",X"11",X"3D",X"8A",X"8A",
		X"5D",X"FB",X"DF",X"DA",X"45",X"5D",X"E2",X"FA",X"A7",X"BB",X"E2",X"BE",X"97",X"2D",X"40",X"FB",
		X"FB",X"5C",X"C7",X"FF",X"97",X"39",X"BF",X"96",X"1D",X"05",X"B7",X"49",X"1D",X"1C",X"53",X"55",
		X"A3",X"B7",X"FC",X"5C",X"FC",X"BB",X"5C",X"00",X"DF",X"15",X"8F",X"7B",X"B9",X"5C",X"9C",X"FF",
		X"1C",X"FA",X"BA",X"01",X"4C",X"BD",X"7A",X"F5",X"34",X"A3",X"6C",X"AB",X"6C",X"49",X"49",X"A1",
		X"71",X"72",X"FC",X"2D",X"72",X"BB",X"75",X"8F",X"35",X"2A",X"B7",X"34",X"E1",X"13",X"E9",X"13",
		X"F1",X"13",X"7F",X"CD",X"35",X"57",X"6E",X"2D",X"02",X"72",X"E3",X"2D",X"8F",X"35",X"19",X"FD",
		X"97",X"A2",X"82",X"FC",X"A3",X"C6",X"FC",X"60",X"9F",X"AE",X"FF",X"E0",X"A3",X"2E",X"FC",X"A2",
		X"99",X"FC",X"FB",X"DB",X"60",X"9F",X"AE",X"BA",X"10",X"ED",X"7A",X"A2",X"46",X"A0",X"37",X"01",
		X"98",X"5F",X"53",X"00",X"8F",X"76",X"FC",X"C1",X"8B",X"B7",X"64",X"E6",X"A3",X"4B",X"FC",X"A3",
		X"0E",X"FC",X"A2",X"99",X"FC",X"4B",X"AF",X"BA",X"FB",X"FB",X"8F",X"FB",X"DC",X"E3",X"9F",X"8B",
		X"B7",X"00",X"8F",X"6B",X"FC",X"A2",X"FF",X"DC",X"60",X"9F",X"AE",X"BB",X"8B",X"8B",X"C7",X"5C",
		X"56",X"EF",X"A3",X"3D",X"B5",X"A2",X"FD",X"FC",X"4B",X"AE",X"DF",X"E2",X"9F",X"5C",X"A6",X"9B",
		X"5C",X"C0",X"8A",X"53",X"A3",X"FD",X"FC",X"A2",X"2F",X"F8",X"60",X"9F",X"AE",X"CA",X"53",X"5C",
		X"D5",X"BB",X"A2",X"FF",X"DC",X"9F",X"9A",X"DC",X"8F",X"9E",X"DC",X"60",X"9F",X"AF",X"FB",X"9F",
		X"BE",X"DC",X"8F",X"FB",X"DC",X"E0",X"E7",X"8B",X"E0",X"79",X"9F",X"CB",X"C1",X"A2",X"3F",X"B5",
		X"69",X"F6",X"68",X"F6",X"DA",X"DA",X"E6",X"D1",X"BA",X"3B",X"BB",X"B6",X"23",X"5C",X"40",X"B2",
		X"A2",X"E2",X"FC",X"60",X"9F",X"AF",X"12",X"5C",X"5C",X"E3",X"5C",X"47",X"92",X"A2",X"A2",X"FC",
		X"4B",X"38",X"BB",X"82",X"53",X"A3",X"B7",X"FC",X"E6",X"A3",X"97",X"FC",X"A3",X"FF",X"DC",X"5C",
		X"61",X"9F",X"53",X"5C",X"D5",X"BB",X"5C",X"CE",X"FB",X"97",X"75",X"B2",X"8F",X"CA",X"B9",X"5C",
		X"9C",X"FF",X"8F",X"A2",X"FC",X"E0",X"4D",X"97",X"69",X"B2",X"8F",X"A5",X"B9",X"60",X"9F",X"AE",
		X"FB",X"97",X"25",X"B2",X"8F",X"27",X"B9",X"5C",X"9C",X"FF",X"0D",X"A2",X"BD",X"B5",X"D9",X"18",
		X"AC",X"FA",X"9F",X"AE",X"BA",X"E0",X"60",X"BB",X"A6",X"CF",X"18",X"A5",X"AF",X"8F",X"FE",X"E0",
		X"17",X"CB",X"C1",X"84",X"A3",X"82",X"FC",X"A3",X"B3",X"FC",X"5C",X"63",X"DB",X"E2",X"9F",X"5C",
		X"A6",X"BA",X"E2",X"BB",X"5C",X"A6",X"BA",X"E2",X"9F",X"A3",X"FD",X"FC",X"19",X"85",X"96",X"A3",
		X"3D",X"B5",X"A2",X"9F",X"FC",X"E6",X"60",X"B7",X"A6",X"BB",X"E2",X"9F",X"A3",X"9F",X"FC",X"5C",
		X"6D",X"FF",X"B6",X"0F",X"8A",X"5D",X"34",X"30",X"05",X"10",X"10",X"8A",X"AA",X"8A",X"AA",X"10",
		X"24",X"15",X"30",X"24",X"8A",X"8A",X"56",X"77",X"34",X"2D",X"15",X"1C",X"05",X"30",X"8A",X"8A",
		X"56",X"77",X"09",X"30",X"77",X"72",X"77",X"34",X"2D",X"15",X"1C",X"05",X"30",X"8A",X"8A",X"53",
		X"5C",X"D5",X"BB",X"A3",X"2F",X"F8",X"8F",X"FF",X"DC",X"E6",X"62",X"97",X"6B",X"FC",X"AE",X"9B",
		X"97",X"2E",X"FC",X"B2",X"4B",X"AE",X"BD",X"A2",X"C6",X"FC",X"60",X"BB",X"AE",X"DF",X"53",X"A3",
		X"E2",X"FC",X"1C",X"E0",X"68",X"9B",X"C1",X"5C",X"61",X"9F",X"E2",X"9B",X"5C",X"A6",X"BA",X"45",
		X"53",X"A3",X"E2",X"FC",X"4D",X"5C",X"D5",X"BB",X"97",X"72",X"92",X"8F",X"C8",X"B9",X"5C",X"9C",
		X"FF",X"0D",X"E0",X"60",X"BB",X"E2",X"A3",X"AE",X"9F",X"C6",X"A3",X"37",X"9D",X"FB",X"67",X"5C",
		X"9E",X"9B",X"05",X"5C",X"A6",X"9B",X"1C",X"4D",X"97",X"5B",X"92",X"8F",X"C8",X"B9",X"5C",X"9C",
		X"FF",X"0D",X"E2",X"9F",X"62",X"E2",X"A3",X"39",X"88",X"92",X"C6",X"A3",X"37",X"9D",X"E2",X"BE",
		X"5C",X"A6",X"BA",X"5C",X"A6",X"9B",X"A2",X"C6",X"FC",X"C6",X"A3",X"C6",X"FC",X"60",X"9F",X"AE",
		X"2B",X"E2",X"9F",X"A3",X"E2",X"FC",X"1C",X"8A",X"71",X"01",X"15",X"0D",X"05",X"77",X"09",X"20",
		X"05",X"30",X"8A",X"AA",X"34",X"2D",X"15",X"1C",X"05",X"30",X"77",X"77",X"8A",X"8A",X"8A",X"65",
		X"01",X"05",X"24",X"77",X"30",X"05",X"15",X"25",X"1C",X"8A",X"AA",X"34",X"2D",X"15",X"1C",X"05",
		X"30",X"77",X"77",X"8A",X"8A",X"53",X"5C",X"D5",X"BB",X"E6",X"A3",X"FF",X"DC",X"5C",X"61",X"9F",
		X"A2",X"A2",X"FC",X"4B",X"AF",X"A2",X"97",X"F5",X"F6",X"8F",X"FA",X"99",X"5C",X"9C",X"FF",X"5C",
		X"CE",X"FB",X"E2",X"AF",X"A3",X"17",X"FC",X"8F",X"B6",X"B9",X"5C",X"E3",X"86",X"FB",X"E6",X"E2",
		X"DB",X"A3",X"9F",X"FC",X"5C",X"6D",X"FF",X"A2",X"A2",X"FC",X"4B",X"AF",X"93",X"5C",X"8F",X"9B",
		X"B7",X"45",X"A2",X"17",X"FC",X"4B",X"AE",X"98",X"71",X"9F",X"CB",X"A3",X"17",X"FC",X"B6",X"51",
		X"53",X"5C",X"D5",X"BB",X"5C",X"CE",X"FB",X"97",X"5E",X"F6",X"8F",X"A8",X"99",X"5C",X"9C",X"FF",
		X"E2",X"D7",X"A3",X"17",X"FC",X"8F",X"B6",X"B9",X"5C",X"E3",X"86",X"FB",X"E6",X"E2",X"DB",X"A3",
		X"9F",X"FC",X"5C",X"6D",X"FF",X"A2",X"BF",X"B5",X"18",X"D8",X"AE",X"D3",X"18",X"D1",X"AE",X"AF",
		X"5C",X"8F",X"9B",X"B7",X"25",X"A2",X"17",X"FC",X"4B",X"AE",X"BE",X"71",X"9F",X"CB",X"A3",X"17",
		X"FC",X"B6",X"31",X"53",X"A3",X"99",X"FC",X"5C",X"63",X"DB",X"E2",X"BA",X"5C",X"A6",X"BA",X"1C",
		X"E2",X"9F",X"B6",X"25",X"8A",X"4D",X"1D",X"29",X"10",X"05",X"30",X"24",X"77",X"11",X"09",X"1D",
		X"29",X"77",X"31",X"05",X"21",X"09",X"30",X"05",X"8A",X"AA",X"77",X"77",X"24",X"1D",X"0D",X"05",
		X"77",X"1D",X"10",X"77",X"04",X"34",X"77",X"24",X"09",X"8A",X"AA",X"77",X"77",X"11",X"09",X"29",
		X"24",X"1D",X"29",X"04",X"05",X"77",X"01",X"15",X"0D",X"05",X"6B",X"8A",X"8A",X"8A",X"71",X"77",
		X"04",X"10",X"05",X"77",X"39",X"09",X"1C",X"10",X"24",X"1D",X"11",X"19",X"77",X"24",X"09",X"77",
		X"10",X"05",X"2D",X"05",X"11",X"24",X"8A",X"AA",X"8A",X"AA",X"8A",X"55",X"10",X"24",X"15",X"30",
		X"24",X"77",X"15",X"24",X"77",X"8A",X"7D",X"6E",X"77",X"77",X"77",X"6A",X"77",X"77",X"8A",X"55",
		X"11",X"09",X"29",X"24",X"1D",X"29",X"04",X"05",X"8A",X"AA",X"2D",X"05",X"20",X"05",X"2D",X"77",
		X"56",X"77",X"77",X"8A",X"7D",X"6E",X"77",X"77",X"77",X"6A",X"77",X"8A",X"55",X"2D",X"15",X"10",
		X"24",X"77",X"01",X"15",X"0D",X"05",X"8A",X"8A",X"93",X"B2",X"4D",X"EB",X"BF",X"C8",X"69",X"3F",
		X"AE",X"9F",X"CF",X"96",X"08",X"0D",X"19",X"29",X"D6",X"4D",X"8B",X"8B",X"E3",X"BF",X"0D",X"1C",
		X"53",X"FA",X"ED",X"01",X"4C",X"B5",X"72",X"4A",X"09",X"8F",X"3C",X"2A",X"6E",X"59",X"58",X"53",
		X"53",X"93",X"53",X"93",X"5F",X"CD",X"34",X"60",X"75",X"08",X"57",X"C3",X"29",X"5C",X"54",X"7D",
		X"75",X"5C",X"8F",X"3C",X"00",X"18",X"E1",X"7D",X"31",X"EA",X"E0",X"4B",X"8A",X"39",X"50",X"D6",
		X"A2",X"E6",X"D8",X"60",X"9B",X"31",X"87",X"F2",X"4D",X"8A",X"8A",X"E3",X"BF",X"5C",X"B9",X"AB",
		X"0D",X"A2",X"BD",X"D8",X"4B",X"3D",X"8B",X"8B",X"C7",X"3D",X"A2",X"3F",X"F8",X"C1",X"8A",X"E3",
		X"3F",X"8A",X"A2",X"E6",X"D8",X"60",X"BB",X"AE",X"CF",X"E3",X"8B",X"8A",X"E3",X"B5",X"8A",X"E3",
		X"FE",X"8A",X"E3",X"DB",X"8A",X"E3",X"2D",X"8A",X"FB",X"AF",X"A2",X"B7",X"FC",X"4B",X"AF",X"BE",
		X"4C",X"D0",X"18",X"D1",X"AE",X"BB",X"FB",X"68",X"A5",X"8A",X"E3",X"FB",X"B6",X"B0",X"A2",X"2B",
		X"F8",X"E6",X"A3",X"2B",X"F8",X"60",X"9A",X"A6",X"9E",X"8B",X"E3",X"BF",X"8A",X"8A",X"8A",X"19",
		X"CE",X"F2",X"E3",X"8B",X"8A",X"E3",X"43",X"8A",X"E3",X"B7",X"8A",X"E3",X"93",X"8A",X"A2",X"B7",
		X"FC",X"4B",X"E2",X"AC",X"FA",X"9B",X"AF",X"AA",X"A2",X"2E",X"F8",X"D9",X"4C",X"D0",X"69",X"DB",
		X"AF",X"9F",X"E6",X"18",X"D1",X"AE",X"BB",X"61",X"24",X"3F",X"60",X"9F",X"21",X"19",X"D6",X"E2",
		X"DF",X"B6",X"FB",X"60",X"FB",X"A6",X"BB",X"E2",X"9F",X"D8",X"DB",X"DB",X"1F",X"DB",X"DB",X"DB",
		X"79",X"25",X"C1",X"8A",X"E3",X"7B",X"8A",X"85",X"8A",X"E3",X"BF",X"9F",X"DB",X"BF",X"9E",X"F1",
		X"8A",X"F0",X"B2",X"60",X"40",X"38",X"04",X"F6",X"60",X"60",X"38",X"2C",X"F6",X"60",X"44",X"4D",
		X"93",X"B2",X"AE",X"9E",X"92",X"8B",X"8B",X"18",X"E1",X"38",X"FD",X"F2",X"B2",X"0D",X"8A",X"C1",
		X"8A",X"8A",X"93",X"B2",X"45",X"7B",X"C1",X"8A",X"93",X"B2",X"7B",X"C1",X"8A",X"8A",X"05",X"7B",
		X"60",X"AE",X"AE",X"8B",X"18",X"C0",X"AF",X"CF",X"C1",X"93",X"8B",X"8B",X"B2",X"7B",X"D9",X"93",
		X"8B",X"B2",X"7B",X"D8",X"93",X"8B",X"8B",X"4D",X"8B",X"81",X"8B",X"A1",X"0D",X"5C",X"B9",X"AB",
		X"1C",X"8A",X"8A",X"E3",X"BF",X"B6",X"61",X"8B",X"E7",X"8A",X"53",X"B6",X"10",X"8B",X"C7",X"8A",
		X"E2",X"EF",X"B6",X"75",X"55",X"4D",X"E0",X"A3",X"E2",X"D8",X"A2",X"B7",X"FC",X"4B",X"AE",X"9E",
		X"5C",X"76",X"82",X"A2",X"C3",X"FC",X"D8",X"B6",X"D8",X"A2",X"E6",X"D8",X"4B",X"AF",X"D9",X"5C",
		X"D2",X"9F",X"A2",X"DE",X"FC",X"D8",X"E2",X"40",X"A3",X"DE",X"FC",X"84",X"CA",X"45",X"A2",X"61",
		X"C7",X"C6",X"C6",X"D8",X"05",X"18",X"C1",X"AE",X"B3",X"D9",X"97",X"24",X"40",X"96",X"E0",X"97",
		X"BE",X"BF",X"96",X"4B",X"A4",X"AF",X"FF",X"18",X"14",X"B6",X"D6",X"69",X"DA",X"AE",X"96",X"18",
		X"15",X"D9",X"69",X"FB",X"AE",X"FB",X"18",X"D1",X"AE",X"FA",X"B6",X"FB",X"18",X"1C",X"18",X"BD",
		X"AE",X"FB",X"18",X"1D",X"B6",X"BB",X"FA",X"3F",X"0D",X"4D",X"A2",X"E6",X"D8",X"4B",X"38",X"7D",
		X"AF",X"97",X"20",X"40",X"96",X"F0",X"8B",X"F1",X"FB",X"DE",X"5C",X"7C",X"8F",X"4B",X"38",X"AC",
		X"D2",X"FB",X"DE",X"5C",X"79",X"8F",X"4B",X"38",X"AC",X"D2",X"8B",X"8B",X"8B",X"8B",X"8B",X"FB",
		X"FF",X"5C",X"7C",X"8F",X"4B",X"AE",X"F7",X"FB",X"FF",X"5C",X"79",X"8F",X"4B",X"AE",X"FE",X"E0",
		X"60",X"3F",X"AE",X"DB",X"E2",X"9F",X"A3",X"2F",X"F8",X"B6",X"C4",X"A2",X"4A",X"F8",X"60",X"3E",
		X"AF",X"E1",X"4D",X"A2",X"E6",X"D8",X"60",X"9F",X"AF",X"9A",X"9F",X"C5",X"BF",X"53",X"5C",X"CA",
		X"DF",X"E2",X"FA",X"B6",X"B8",X"60",X"BB",X"AF",X"A7",X"A2",X"0B",X"F8",X"E6",X"A3",X"0B",X"F8",
		X"60",X"BA",X"AF",X"B2",X"E2",X"D7",X"5C",X"A6",X"BA",X"A2",X"FF",X"DC",X"60",X"9F",X"9F",X"6B",
		X"FC",X"AE",X"9B",X"9F",X"2E",X"FC",X"BA",X"E6",X"BB",X"5C",X"1F",X"DF",X"E2",X"B7",X"D9",X"FA",
		X"BF",X"53",X"5C",X"CA",X"DF",X"E2",X"DE",X"B6",X"F3",X"9F",X"BF",X"BB",X"53",X"5C",X"CA",X"DF",
		X"A2",X"DD",X"D8",X"68",X"9F",X"4B",X"A3",X"DD",X"D8",X"E2",X"FE",X"AE",X"BB",X"E2",X"96",X"5C",
		X"A6",X"BA",X"5C",X"E6",X"EA",X"0D",X"FA",X"3D",X"07",X"C1",X"5C",X"31",X"EA",X"1D",X"1D",X"1D",
		X"9F",X"00",X"40",X"9E",X"93",X"19",X"9B",X"F2",X"0D",X"4D",X"5C",X"74",X"8F",X"A2",X"E6",X"D8",
		X"60",X"9F",X"38",X"5E",X"8F",X"0D",X"4D",X"E0",X"60",X"37",X"39",X"40",X"D2",X"84",X"60",X"37",
		X"38",X"5E",X"8F",X"FB",X"DF",X"5C",X"E0",X"DB",X"8B",X"8B",X"E8",X"EB",X"DC",X"E0",X"E3",X"BF",
		X"69",X"D2",X"C6",X"8B",X"F9",X"0D",X"4D",X"97",X"04",X"40",X"96",X"D1",X"E0",X"D0",X"DB",X"DB",
		X"1B",X"4C",X"FD",X"D0",X"EB",X"BF",X"AC",X"8E",X"8E",X"A0",X"F3",X"40",X"96",X"97",X"9A",X"FD",
		X"96",X"5D",X"4D",X"D0",X"DB",X"1B",X"F3",X"BF",X"D0",X"8F",X"88",X"EF",X"96",X"F9",X"F3",X"BF",
		X"B4",X"8B",X"F8",X"0D",X"4D",X"A2",X"2D",X"DC",X"C1",X"8A",X"B7",X"64",X"55",X"97",X"2D",X"40",
		X"96",X"15",X"96",X"99",X"DE",X"AF",X"05",X"0D",X"97",X"BF",X"64",X"96",X"08",X"8F",X"36",X"DC",
		X"4D",X"E0",X"4B",X"AE",X"F3",X"8B",X"8B",X"E0",X"02",X"AF",X"DF",X"8B",X"E0",X"22",X"AE",X"DB",
		X"0D",X"8B",X"8B",X"8B",X"8B",X"B6",X"0C",X"8A",X"8A",X"E3",X"40",X"0D",X"1D",X"0D",X"4D",X"97",
		X"24",X"40",X"96",X"E0",X"4B",X"39",X"16",X"AF",X"8B",X"84",X"69",X"2F",X"60",X"2F",X"AF",X"CF",
		X"F9",X"A2",X"2E",X"F8",X"37",X"60",X"40",X"AE",X"FB",X"60",X"9F",X"18",X"1D",X"AF",X"F7",X"8B",
		X"F9",X"A2",X"0E",X"F8",X"37",X"18",X"C0",X"AE",X"BB",X"4C",X"FD",X"D9",X"A2",X"5F",X"F8",X"26",
		X"31",X"5E",X"8F",X"FA",X"37",X"84",X"60",X"37",X"39",X"7D",X"AF",X"0D",X"4D",X"97",X"20",X"40",
		X"96",X"F9",X"8A",X"E0",X"C6",X"D0",X"DB",X"1B",X"DB",X"1B",X"DB",X"F3",X"BF",X"D0",X"8F",X"B7",
		X"DC",X"96",X"8B",X"E0",X"8B",X"4B",X"AE",X"9D",X"37",X"18",X"C0",X"AE",X"BB",X"4C",X"FD",X"60",
		X"9E",X"A7",X"48",X"8A",X"F1",X"8A",X"E0",X"18",X"C0",X"AF",X"EA",X"4B",X"AE",X"8A",X"AB",X"F9",
		X"D8",X"D4",X"55",X"C6",X"D0",X"DB",X"1B",X"F3",X"BF",X"D0",X"8F",X"A8",X"EF",X"96",X"E0",X"15",
		X"3B",X"37",X"18",X"C0",X"AE",X"BB",X"4C",X"FD",X"60",X"FF",X"A7",X"DE",X"AA",X"F9",X"D8",X"18",
		X"60",X"0D",X"4D",X"8B",X"8B",X"81",X"19",X"5E",X"8F",X"0D",X"4D",X"E0",X"D8",X"69",X"7B",X"60",
		X"7B",X"AF",X"F7",X"A2",X"B7",X"FC",X"4B",X"AF",X"A2",X"4C",X"D0",X"69",X"C2",X"60",X"9B",X"A7",
		X"A3",X"84",X"68",X"9F",X"D8",X"B6",X"EE",X"4C",X"D0",X"69",X"C2",X"60",X"AF",X"FA",X"7B",X"A6",
		X"AB",X"FE",X"B6",X"D2",X"0D",X"4D",X"A2",X"E6",X"D8",X"4B",X"AF",X"FA",X"97",X"24",X"40",X"96",
		X"E0",X"4B",X"AF",X"FB",X"84",X"60",X"3E",X"38",X"5E",X"8F",X"0D",X"4D",X"84",X"69",X"7B",X"60",
		X"7B",X"AF",X"B8",X"97",X"24",X"40",X"96",X"E0",X"4B",X"39",X"5E",X"8F",X"8B",X"8B",X"E0",X"79",
		X"BE",X"D9",X"8A",X"E0",X"18",X"9D",X"AF",X"FF",X"C6",X"38",X"B2",X"8F",X"C6",X"D0",X"DB",X"1B",
		X"DB",X"F3",X"BF",X"D0",X"8F",X"B4",X"DC",X"96",X"E0",X"8B",X"4B",X"AE",X"DE",X"37",X"18",X"C0",
		X"AE",X"BB",X"4C",X"FD",X"60",X"DB",X"A7",X"25",X"B6",X"81",X"A2",X"E6",X"D8",X"4B",X"AE",X"88",
		X"4C",X"D0",X"69",X"C2",X"60",X"AF",X"FA",X"7F",X"A6",X"F7",X"FE",X"B6",X"97",X"0D",X"4D",X"97",
		X"24",X"40",X"96",X"84",X"69",X"7B",X"60",X"7F",X"AF",X"95",X"E0",X"4B",X"AF",X"A2",X"0D",X"4D",
		X"97",X"20",X"40",X"96",X"E0",X"79",X"BE",X"18",X"9D",X"AE",X"BB",X"71",X"B7",X"D9",X"8A",X"E0",
		X"C6",X"D0",X"DB",X"1B",X"DB",X"F3",X"BF",X"D0",X"8F",X"A4",X"DC",X"96",X"E0",X"8B",X"4B",X"AE",
		X"EE",X"37",X"18",X"C0",X"AE",X"BB",X"4C",X"FD",X"60",X"FF",X"A7",X"25",X"A2",X"E6",X"D8",X"4B",
		X"AE",X"96",X"84",X"68",X"9F",X"D8",X"B6",X"D7",X"A2",X"E6",X"D8",X"4B",X"AF",X"DE",X"E0",X"60",
		X"FF",X"FA",X"7B",X"AE",X"BE",X"60",X"EF",X"FA",X"5B",X"AE",X"BB",X"FA",X"3F",X"0D",X"84",X"A3",
		X"C2",X"D8",X"A2",X"E2",X"D8",X"06",X"15",X"B2",X"38",X"44",X"D6",X"85",X"4D",X"A2",X"E6",X"D8",
		X"DB",X"F3",X"BF",X"D0",X"8F",X"7E",X"AB",X"96",X"F0",X"8B",X"F1",X"84",X"5C",X"90",X"AB",X"DB",
		X"EB",X"BF",X"C8",X"96",X"F0",X"8B",X"F1",X"5C",X"7F",X"AB",X"0D",X"8A",X"A1",X"8A",X"81",X"0D",
		X"92",X"E2",X"44",X"19",X"09",X"D6",X"A2",X"2A",X"F8",X"33",X"B6",X"FF",X"A2",X"0E",X"F8",X"13",
		X"18",X"C0",X"AE",X"BB",X"4C",X"FD",X"26",X"E2",X"BF",X"35",X"E6",X"1C",X"A2",X"B7",X"FC",X"4B",
		X"3D",X"F8",X"8B",X"C7",X"3D",X"A2",X"3F",X"F8",X"D0",X"4C",X"D0",X"69",X"C2",X"60",X"B7",X"A7",
		X"9F",X"F6",X"81",X"8A",X"A2",X"E6",X"D8",X"60",X"9F",X"AE",X"FB",X"60",X"BB",X"AE",X"A3",X"B6",
		X"AB",X"A2",X"0E",X"F8",X"D9",X"A2",X"67",X"F8",X"97",X"BF",X"BF",X"FA",X"7F",X"26",X"A6",X"BB",
		X"FE",X"F7",X"A2",X"2A",X"F8",X"D9",X"A2",X"47",X"F8",X"26",X"A7",X"9F",X"F6",X"80",X"2A",X"3D",
		X"18",X"1C",X"1C",X"FA",X"2F",X"4C",X"D0",X"69",X"FE",X"3D",X"FA",X"37",X"4C",X"D0",X"69",X"FB",
		X"3D",X"E0",X"69",X"9F",X"FA",X"7B",X"07",X"D8",X"4C",X"D0",X"69",X"DB",X"3D",X"84",X"68",X"9F",
		X"D8",X"1C",X"4D",X"A2",X"C6",X"D8",X"DB",X"DB",X"D0",X"F3",X"BF",X"8F",X"7B",X"F8",X"96",X"15",
		X"B2",X"C1",X"8B",X"92",X"B2",X"C1",X"8B",X"A5",X"8B",X"85",X"1C",X"5D",X"FB",X"9E",X"18",X"C1",
		X"AF",X"B6",X"DF",X"18",X"C8",X"AF",X"F3",X"DF",X"DF",X"18",X"C9",X"AF",X"DE",X"DF",X"18",X"D0",
		X"AF",X"BE",X"DF",X"18",X"D1",X"AE",X"9B",X"69",X"9B",X"D9",X"A4",X"1D",X"1C",X"18",X"D9",X"AF",
		X"04",X"DF",X"B6",X"61",X"E2",X"40",X"22",X"3D",X"B6",X"60",X"40",X"40",X"72",X"AB",X"DE",X"8B",
		X"AD",X"8B",X"62",X"8B",X"62",X"8B",X"62",X"8B",X"62",X"8B",X"62",X"8B",X"62",X"8B",X"07",X"AB",
		X"39",X"AB",X"11",X"AB",X"50",X"AB",X"08",X"AB",X"41",X"AB",X"3A",X"AB",X"3A",X"AB",X"3A",X"3A",
		X"AB",X"F9",X"BF",X"BB",X"BF",X"BF",X"B8",X"BF",X"BB",X"60",X"BF",X"F8",X"BF",X"BB",X"44",X"BF",
		X"60",X"25",X"FD",X"BF",X"60",X"BF",X"BF",X"BC",X"BF",X"60",X"BB",X"BF",X"FC",X"BF",X"60",X"9B",
		X"BF",X"60",X"25",X"B5",X"64",X"BF",X"BF",X"BF",X"FD",X"64",X"BF",X"BF",X"BF",X"60",X"45",X"B5",
		X"FF",X"BF",X"BF",X"BF",X"FD",X"FF",X"BF",X"BF",X"BF",X"60",X"45",X"FD",X"BF",X"BF",X"BF",X"BF",
		X"F9",X"BF",X"BF",X"BF",X"BF",X"60",X"45",X"F5",X"BF",X"BF",X"BF",X"BF",X"F9",X"BF",X"BF",X"BF",
		X"BF",X"F1",X"BF",X"BF",X"BF",X"BF",X"FD",X"BF",X"BF",X"BF",X"BF",X"60",X"08",X"AF",X"8B",X"EE",
		X"8B",X"A6",X"8B",X"FD",X"8B",X"B5",X"8B",X"3A",X"AB",X"3A",X"AB",X"3A",X"AB",X"3A",X"3A",X"AB",
		X"FB",X"FF",X"FF",X"BF",X"BF",X"BA",X"FF",X"FF",X"BF",X"BF",X"60",X"45",X"FF",X"64",X"64",X"BF",
		X"BF",X"BE",X"64",X"64",X"BF",X"BF",X"60",X"45",X"FB",X"64",X"FF",X"BF",X"BF",X"BA",X"64",X"FF",
		X"BF",X"BF",X"60",X"45",X"FF",X"FF",X"64",X"BF",X"BF",X"BE",X"FF",X"64",X"BF",X"BF",X"60",X"45",
		X"FE",X"BF",X"BF",X"BF",X"BF",X"FA",X"BF",X"BF",X"BF",X"BF",X"60",X"45",X"00",X"19",X"1A",X"CF",
		X"81",X"8B",X"7F",X"8B",X"57",X"8B",X"6B",X"8B",X"43",X"8B",X"3A",X"AB",X"3A",X"AB",X"3A",X"AB",
		X"3A",X"3A",X"AB",X"B3",X"BF",X"BB",X"BF",X"BE",X"F3",X"BF",X"BB",X"BF",X"9E",X"B2",X"BF",X"FF",
		X"BF",X"BA",X"60",X"25",X"B7",X"BF",X"60",X"BF",X"BE",X"F7",X"BF",X"60",X"BF",X"DB",X"B6",X"BF",
		X"64",X"BF",X"9E",X"60",X"25",X"B7",X"64",X"BF",X"BF",X"FB",X"F7",X"64",X"BF",X"BF",X"DB",X"B6",
		X"64",X"BF",X"BF",X"BE",X"60",X"45",X"B7",X"FF",X"BF",X"BF",X"BE",X"F7",X"FF",X"BF",X"BF",X"DB",
		X"B6",X"FF",X"BF",X"BF",X"FB",X"60",X"45",X"B7",X"BF",X"BF",X"BF",X"BE",X"60",X"20",X"31",X"8B",
		X"2C",X"8B",X"60",X"8B",X"BA",X"EF",X"89",X"EF",X"3A",X"AB",X"F3",X"EF",X"CB",X"EF",X"F9",X"EF",
		X"3A",X"AB",X"B0",X"BF",X"9B",X"BF",X"BF",X"F0",X"BF",X"9B",X"BF",X"BF",X"A9",X"BF",X"BB",X"BF",
		X"BF",X"E9",X"BF",X"BB",X"BF",X"BF",X"60",X"08",X"B4",X"BF",X"44",X"BF",X"BF",X"F4",X"BF",X"44",
		X"BF",X"BF",X"AD",X"BF",X"60",X"BF",X"BF",X"ED",X"BF",X"60",X"BF",X"BF",X"60",X"08",X"B4",X"64",
		X"BF",X"BF",X"BF",X"AC",X"64",X"BF",X"BF",X"BF",X"60",X"45",X"B4",X"FF",X"BF",X"BF",X"BF",X"AC",
		X"FF",X"BF",X"BF",X"BF",X"60",X"45",X"B4",X"BF",X"BF",X"BF",X"BF",X"EC",X"BF",X"BF",X"BF",X"BF",
		X"A5",X"BF",X"BF",X"BF",X"BF",X"60",X"25",X"E5",X"64",X"BF",X"BF",X"BF",X"44",X"E5",X"20",X"BF",
		X"BF",X"BF",X"44",X"E5",X"24",X"BF",X"BF",X"BF",X"44",X"E5",X"61",X"BF",X"BF",X"BF",X"44",X"E5",
		X"65",X"BF",X"BF",X"BF",X"60",X"F2",X"A4",X"FF",X"BF",X"BF",X"BF",X"44",X"A4",X"FB",X"BF",X"BF",
		X"BF",X"44",X"A4",X"BE",X"BF",X"BF",X"BF",X"44",X"A4",X"BA",X"BF",X"BF",X"BF",X"44",X"A4",X"FE",
		X"BF",X"BF",X"BF",X"B4",X"BF",X"BF",X"BF",X"BF",X"60",X"20",X"BF",X"BB",X"BB",X"BF",X"BB",X"BB",
		X"24",X"BB",X"FF",X"FF",X"9F",X"9F",X"64",X"9B",X"9B",X"BF",X"9B",X"BB",X"BF",X"BB",X"BB",X"BF",
		X"9B",X"BB",X"BF",X"BB",X"BB",X"BF",X"9B",X"BB",X"BF",X"9B",X"BB",X"BF",X"9B",X"BB",X"BF",X"BB",
		X"BB",X"64",X"FF",X"9B",X"BF",X"FF",X"BB",X"BF",X"FF",X"BB",X"BF",X"9B",X"BB",X"53",X"5C",X"D5",
		X"BB",X"5C",X"D0",X"BB",X"FB",X"F2",X"5C",X"9E",X"9B",X"01",X"10",X"C8",X"41",X"DF",X"69",X"A8",
		X"DD",X"F9",X"C0",X"83",X"DB",X"F5",X"26",X"F3",X"0D",X"A8",X"F3",X"72",X"A8",X"E6",X"DB",X"83",
		X"E2",X"CD",X"DB",X"83",X"DF",X"26",X"C6",X"FB",X"F6",X"AC",X"0E",X"B4",X"00",X"A2",X"FF",X"DC",
		X"60",X"9F",X"9F",X"BD",X"FC",X"97",X"0B",X"FC",X"8F",X"FB",X"DC",X"AE",X"9E",X"9F",X"9D",X"FC",
		X"97",X"6F",X"FC",X"8F",X"9E",X"DC",X"B2",X"A3",X"4F",X"FC",X"BA",X"A3",X"B9",X"FC",X"4B",X"AF",
		X"97",X"9F",X"CC",X"F8",X"A2",X"FF",X"DC",X"60",X"9F",X"AE",X"9B",X"9F",X"E5",X"F8",X"BA",X"A3",
		X"2B",X"F8",X"E0",X"60",X"F7",X"AF",X"97",X"A2",X"B7",X"FC",X"4B",X"E0",X"AF",X"BA",X"A2",X"4F",
		X"FC",X"E6",X"A3",X"4F",X"FC",X"E2",X"9F",X"C1",X"97",X"5C",X"CA",X"C6",X"DB",X"EB",X"BF",X"C8",
		X"96",X"E0",X"8B",X"E9",X"C8",X"5C",X"E8",X"8A",X"A3",X"2D",X"DC",X"79",X"F6",X"A3",X"50",X"DC",
		X"4D",X"5C",X"23",X"BB",X"19",X"3D",X"CA",X"EF",X"B6",X"2D",X"40",X"CD",X"99",X"EF",X"F7",X"2D",
		X"40",X"EF",X"99",X"EF",X"B7",X"2D",X"40",X"09",X"B9",X"EF",X"FE",X"2D",X"40",X"2B",X"B9",X"EF",
		X"BA",X"2D",X"40",X"1F",X"B9",X"EF",X"BE",X"2D",X"40",X"AD",X"B9",X"AB",X"FF",X"42",X"40",X"4F",
		X"99",X"EB",X"FF",X"C2",X"BF",X"DD",X"BD",X"8B",X"FF",X"42",X"40",X"5F",X"99",X"CF",X"FF",X"C2",
		X"BF",X"CD",X"BD",X"EE",X"BB",X"50",X"40",X"0F",X"B9",X"CA",X"BB",X"D2",X"BF",X"9D",X"9D",X"8A",
		X"58",X"4B",X"67",X"67",X"67",X"67",X"67",X"67",X"6F",X"8A",X"8A",X"A2",X"BA",X"FC",X"D9",X"A2",
		X"9A",X"FC",X"97",X"2D",X"40",X"8F",X"7B",X"99",X"5D",X"45",X"01",X"10",X"3C",X"7A",X"82",X"46",
		X"4E",X"49",X"49",X"01",X"98",X"8D",X"00",X"05",X"5C",X"C7",X"FF",X"9F",X"DD",X"9B",X"9E",X"1D",
		X"B7",X"69",X"E2",X"AA",X"A3",X"42",X"99",X"E2",X"8A",X"A3",X"D0",X"BD",X"E2",X"82",X"97",X"2D",
		X"40",X"8F",X"52",X"99",X"FB",X"B2",X"5C",X"C7",X"FF",X"8F",X"E3",X"CF",X"FB",X"FE",X"5D",X"8B",
		X"E0",X"8B",X"F9",X"8B",X"F0",X"8B",X"F1",X"8B",X"F8",X"8B",X"4D",X"E9",X"8C",X"5D",X"4D",X"5C",
		X"C7",X"FF",X"0D",X"9F",X"BF",X"FF",X"9E",X"1D",X"E2",X"92",X"5C",X"C7",X"FF",X"0D",X"1D",X"B7",
		X"54",X"97",X"C0",X"CF",X"8F",X"6C",X"99",X"5C",X"99",X"FF",X"E2",X"EF",X"A3",X"78",X"99",X"A3",
		X"15",X"99",X"E2",X"97",X"A3",X"78",X"D9",X"A3",X"15",X"D9",X"0D",X"8B",X"FB",X"DF",X"97",X"BA",
		X"D8",X"4C",X"91",X"80",X"F8",X"97",X"36",X"DC",X"4C",X"91",X"73",X"DC",X"97",X"3C",X"F8",X"4C",
		X"91",X"14",X"DC",X"A2",X"FF",X"DC",X"60",X"9F",X"97",X"E8",X"F8",X"AE",X"9B",X"97",X"C5",X"F8",
		X"4C",X"91",X"10",X"DC",X"97",X"2A",X"99",X"5D",X"55",X"E2",X"68",X"A3",X"DE",X"DC",X"A4",X"A3",
		X"FE",X"DC",X"4D",X"C6",X"D8",X"DB",X"1F",X"DB",X"45",X"FB",X"BF",X"D8",X"8F",X"B4",X"DC",X"9E",
		X"AB",X"F1",X"DC",X"8F",X"A4",X"DC",X"9E",X"AB",X"E1",X"DC",X"A2",X"FE",X"DC",X"C6",X"D8",X"05",
		X"1F",X"DB",X"D8",X"A2",X"FF",X"DC",X"60",X"9F",X"8F",X"0D",X"DC",X"AE",X"9B",X"8F",X"CB",X"F8",
		X"9E",X"AB",X"54",X"DC",X"8F",X"B7",X"DC",X"9E",X"AB",X"FA",X"DC",X"0D",X"5C",X"E8",X"8A",X"8B",
		X"DB",X"DB",X"DB",X"DB",X"FB",X"FF",X"5C",X"52",X"CB",X"5C",X"E8",X"8A",X"8B",X"FB",X"BE",X"5C",
		X"52",X"CB",X"5C",X"E8",X"8A",X"8B",X"FB",X"BE",X"5C",X"52",X"CB",X"5C",X"E8",X"8A",X"8B",X"FB",
		X"BE",X"5C",X"52",X"CB",X"4D",X"53",X"AA",X"F1",X"DC",X"C1",X"AA",X"E1",X"DC",X"C1",X"AA",X"FA",
		X"DC",X"8B",X"C1",X"0D",X"15",X"93",X"93",X"93",X"93",X"93",X"1D",X"DF",X"39",X"C3",X"EB",X"AA",
		X"73",X"DC",X"E3",X"BF",X"8F",X"4B",X"F8",X"53",X"C1",X"8B",X"E6",X"C1",X"8B",X"E3",X"69",X"8B",
		X"E3",X"B6",X"8B",X"E3",X"BA",X"8B",X"E3",X"FF",X"8B",X"E3",X"08",X"8B",X"E3",X"AB",X"8B",X"E3",
		X"3F",X"A2",X"FF",X"DC",X"60",X"9F",X"97",X"0B",X"FC",X"8F",X"BE",X"DC",X"AE",X"FB",X"97",X"6F",
		X"FC",X"8F",X"9A",X"DC",X"A2",X"4F",X"FC",X"B3",X"E0",X"60",X"B7",X"A6",X"BA",X"A2",X"B7",X"FC",
		X"4B",X"E0",X"AF",X"9B",X"E2",X"DA",X"C1",X"97",X"24",X"C7",X"C6",X"DB",X"EB",X"BF",X"C8",X"96",
		X"E0",X"8B",X"E9",X"C8",X"A2",X"4F",X"FC",X"4B",X"E0",X"AE",X"9F",X"53",X"9F",X"C4",X"F8",X"BB",
		X"8B",X"E0",X"9B",X"BB",X"9B",X"BB",X"8B",X"E0",X"9B",X"BB",X"8B",X"E0",X"9B",X"BB",X"A3",X"02",
		X"F8",X"8B",X"E0",X"9B",X"BB",X"8B",X"E0",X"9B",X"BB",X"A3",X"79",X"F8",X"8B",X"E0",X"9B",X"BB",
		X"8B",X"E0",X"9B",X"BB",X"A2",X"4F",X"FC",X"4B",X"AE",X"FF",X"8F",X"E0",X"F8",X"C7",X"A2",X"B7",
		X"FC",X"4B",X"AF",X"A2",X"E2",X"9F",X"A3",X"BF",X"FC",X"5C",X"F7",X"DF",X"5C",X"3E",X"DF",X"5C",
		X"11",X"DF",X"A2",X"82",X"FC",X"60",X"BB",X"AF",X"9E",X"5C",X"F6",X"DF",X"5C",X"77",X"DF",X"5C",
		X"70",X"DF",X"E2",X"FF",X"A3",X"BF",X"FC",X"5C",X"7C",X"DF",X"A2",X"4A",X"FC",X"4B",X"AF",X"FA",
		X"8F",X"9D",X"D8",X"E3",X"BB",X"8B",X"E3",X"B5",X"8B",X"E3",X"BF",X"5C",X"24",X"FB",X"1C",X"AA",
		X"14",X"DC",X"55",X"97",X"BE",X"BF",X"96",X"E3",X"BF",X"8B",X"8B",X"8B",X"15",X"B6",X"C8",X"5D",
		X"55",X"DB",X"31",X"15",X"AE",X"45",X"5C",X"E8",X"8A",X"8B",X"4D",X"18",X"C0",X"AE",X"89",X"18",
		X"42",X"45",X"A2",X"B9",X"FC",X"4B",X"AF",X"DA",X"AA",X"10",X"DC",X"E0",X"8B",X"AB",X"10",X"DC",
		X"18",X"C1",X"AF",X"18",X"4B",X"AE",X"3C",X"8F",X"72",X"F8",X"E7",X"8F",X"52",X"F8",X"E7",X"AA",
		X"14",X"DC",X"A2",X"FE",X"DC",X"D8",X"DB",X"DB",X"1F",X"DB",X"DB",X"DB",X"79",X"25",X"D9",X"E3",
		X"BF",X"8B",X"85",X"8B",X"A2",X"DE",X"DC",X"C1",X"8B",X"A5",X"8B",X"A2",X"2D",X"DC",X"60",X"9B",
		X"FB",X"D3",X"AE",X"BE",X"60",X"BB",X"FB",X"DE",X"AE",X"BB",X"FB",X"B7",X"A5",X"8B",X"E3",X"B6",
		X"8B",X"E3",X"89",X"8B",X"E3",X"EF",X"8B",X"E3",X"3F",X"8B",X"E3",X"BA",X"8B",X"8B",X"AB",X"14",
		X"DC",X"05",X"18",X"C1",X"AE",X"9A",X"18",X"43",X"AA",X"E1",X"DC",X"5C",X"04",X"AE",X"AB",X"E1",
		X"DC",X"4B",X"38",X"58",X"AE",X"60",X"F2",X"AF",X"93",X"45",X"93",X"A2",X"FE",X"DC",X"60",X"9F",
		X"E2",X"BE",X"AF",X"BB",X"E2",X"82",X"B3",X"92",X"05",X"19",X"42",X"AE",X"60",X"D2",X"AF",X"D2",
		X"D9",X"8F",X"0F",X"F8",X"E7",X"AA",X"80",X"F8",X"A2",X"FE",X"DC",X"C1",X"8B",X"A2",X"DE",X"DC",
		X"C1",X"8B",X"81",X"8B",X"A1",X"8B",X"E3",X"9F",X"8B",X"AB",X"80",X"F8",X"A4",X"B6",X"AD",X"60",
		X"B3",X"AF",X"9A",X"AA",X"F1",X"DC",X"5C",X"04",X"AE",X"AB",X"F1",X"DC",X"B6",X"95",X"FA",X"BF",
		X"60",X"B3",X"A7",X"BB",X"18",X"1D",X"60",X"9A",X"A6",X"FB",X"60",X"D7",X"A7",X"BB",X"18",X"1C",
		X"18",X"9D",X"AE",X"D6",X"D9",X"A2",X"B9",X"FC",X"4B",X"AF",X"FE",X"AA",X"54",X"DC",X"E0",X"8B",
		X"8B",X"AB",X"54",X"DC",X"4B",X"AE",X"B1",X"A4",X"AA",X"FA",X"DC",X"5C",X"41",X"AE",X"AB",X"FA",
		X"DC",X"18",X"9C",X"AE",X"B2",X"45",X"71",X"9A",X"FB",X"BF",X"D8",X"8F",X"9F",X"8E",X"9E",X"F9",
		X"AA",X"73",X"DC",X"A5",X"8B",X"C1",X"8B",X"81",X"8B",X"A1",X"8B",X"AB",X"73",X"DC",X"05",X"8F",
		X"BE",X"8E",X"C6",X"DB",X"FB",X"BF",X"D8",X"9E",X"E0",X"8B",X"E9",X"C8",X"5C",X"0B",X"FF",X"0D",
		X"05",X"15",X"4D",X"8F",X"2D",X"40",X"96",X"08",X"0D",X"45",X"A2",X"DE",X"DC",X"71",X"BE",X"A3",
		X"DE",X"DC",X"05",X"1D",X"DF",X"39",X"52",X"CB",X"1C",X"AA",X"FA",X"DC",X"E3",X"BF",X"8B",X"E3",
		X"40",X"8B",X"AB",X"FA",X"DC",X"B6",X"34",X"C1",X"8B",X"45",X"A2",X"DE",X"DC",X"C1",X"8B",X"05",
		X"1C",X"D5",X"40",X"D5",X"D5",X"9B",X"B8",X"97",X"F9",X"8E",X"B5",X"8E",X"B0",X"8E",X"EC",X"8E",
		X"A5",X"8E",X"7F",X"8E",X"33",X"8E",X"76",X"8E",X"2A",X"8E",X"67",X"8E",X"39",X"8E",X"35",X"8E",
		X"70",X"8E",X"2C",X"8E",X"BB",X"AA",X"F7",X"AA",X"EB",X"AA",X"E7",X"AA",X"F0",X"AA",X"AC",X"AA",
		X"A1",X"AA",X"3E",X"AA",X"72",X"AA",X"2A",X"AA",X"63",X"AA",X"39",X"AA",X"78",X"AA",X"30",X"AA",
		X"69",X"AA",X"64",X"AA",X"BE",X"8A",X"BB",X"BB",X"7A",X"9A",X"7E",X"9A",X"5A",X"9A",X"5E",X"9A",
		X"BB",X"BB",X"3A",X"9A",X"3E",X"FE",X"1A",X"9A",X"1E",X"FE",X"BB",X"FF",X"7F",X"9A",X"3F",X"FE",
		X"5F",X"9A",X"1F",X"FE",X"7B",X"9A",X"3B",X"FE",X"5B",X"9A",X"1B",X"FE",X"9F",X"9F",X"47",X"9A",
		X"9B",X"9B",X"65",X"97",X"05",X"97",X"BF",X"BF",X"BF",X"BF",X"21",X"97",X"25",X"B2",X"45",X"97",
		X"01",X"97",X"BF",X"BF",X"9B",X"BB",X"2E",X"FF",X"6B",X"F2",X"6F",X"9E",X"0E",X"BE",X"4B",X"FA",
		X"4F",X"9E",X"BB",X"BB",X"33",X"92",X"37",X"DF",X"13",X"92",X"17",X"DF",X"9B",X"BB",X"2B",X"FA",
		X"2F",X"FA",X"72",X"FA",X"0B",X"FA",X"0F",X"FA",X"52",X"FA",X"BB",X"BB",X"73",X"97",X"77",X"D6",
		X"53",X"97",X"57",X"D6",X"9B",X"BB",X"76",X"FA",X"32",X"97",X"36",X"97",X"56",X"FA",X"12",X"97",
		X"16",X"97",X"9B",X"BB",X"7C",X"97",X"38",X"B2",X"3C",X"D3",X"5C",X"97",X"18",X"B2",X"1C",X"D3",
		X"9B",X"BB",X"7D",X"FE",X"39",X"96",X"3D",X"96",X"5D",X"FE",X"19",X"96",X"1D",X"96",X"BB",X"BB",
		X"31",X"F7",X"35",X"DE",X"11",X"F7",X"15",X"DE",X"FF",X"9B",X"0C",X"93",X"69",X"DA",X"09",X"DA",
		X"2D",X"DA",X"28",X"F7",X"49",X"F6",X"6D",X"B3",X"0D",X"DA",X"08",X"93",X"2C",X"B3",X"4D",X"B3",
		X"29",X"B3",X"FF",X"BB",X"BF",X"BF",X"BF",X"BF",X"30",X"B6",X"34",X"B6",X"BF",X"BF",X"BF",X"BF",
		X"10",X"B6",X"14",X"B6",X"FF",X"BB",X"62",X"DB",X"66",X"F6",X"22",X"D3",X"26",X"D3",X"42",X"DB",
		X"46",X"F6",X"02",X"D3",X"06",X"D3",X"9B",X"BB",X"6A",X"FF",X"6E",X"FF",X"2A",X"FF",X"4A",X"FF",
		X"4E",X"FF",X"0A",X"FF",X"DF",X"FF",X"F7",X"D7",X"93",X"97",X"B3",X"97",X"97",X"97",X"B7",X"BF",
		X"D3",X"D7",X"F3",X"D7",X"D7",X"9A",X"D7",X"9A",X"D7",X"9A",X"D3",X"D7",X"F2",X"D7",X"D6",X"9A",
		X"D6",X"9A",X"D6",X"9A",X"F6",X"D7",X"92",X"97",X"B2",X"97",X"96",X"97",X"B6",X"BF",X"FF",X"9F",
		X"AF",X"BF",X"AF",X"BF",X"A0",X"BF",X"A1",X"FB",X"FF",X"9F",X"AF",X"BF",X"AF",X"BF",X"C4",X"BF",
		X"C5",X"FB",X"DF",X"BB",X"BB",X"BF",X"BB",X"BF",X"BB",X"BF",X"A4",X"BF",X"A5",X"BF",X"AF",X"BF",
		X"AF",X"BF",X"AF",X"BF",X"AF",X"BF",X"85",X"BF",X"DF",X"BB",X"AF",X"BF",X"AF",X"BF",X"AF",X"BF",
		X"AF",X"BF",X"E1",X"BF",X"9B",X"BF",X"9B",X"BF",X"9B",X"BF",X"C0",X"BF",X"C1",X"BF",X"DF",X"9F",
		X"E5",X"BF",X"E5",X"BF",X"E5",X"BF",X"E5",X"BF",X"E4",X"BF",X"DF",X"9F",X"81",X"BF",X"81",X"BF",
		X"81",X"BF",X"81",X"BF",X"80",X"BF",X"DF",X"9F",X"9B",X"BF",X"9B",X"BF",X"9B",X"BF",X"9B",X"BF",
		X"9A",X"BF",X"DF",X"9F",X"BB",X"BF",X"BB",X"BF",X"BB",X"BF",X"BB",X"BF",X"BA",X"BF",X"DF",X"9F",
		X"E5",X"BF",X"E5",X"BF",X"E5",X"BF",X"E5",X"BF",X"E5",X"BF",X"DF",X"9F",X"81",X"BF",X"81",X"BF",
		X"81",X"BF",X"81",X"BF",X"81",X"BF",X"DF",X"BB",X"9B",X"BF",X"9B",X"BF",X"9B",X"BF",X"9B",X"BF",
		X"9A",X"BF",X"BB",X"BF",X"BB",X"BF",X"BB",X"BF",X"BB",X"BF",X"BA",X"BF",X"DF",X"9F",X"BF",X"BF",
		X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BE",X"BF",X"DF",X"BB",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",
		X"ED",X"F3",X"BE",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"BF",X"CD",X"F3",X"CC",X"BF",X"BF",X"BF",
		X"BF",X"BF",X"E8",X"F3",X"E9",X"F3",X"BE",X"BF",X"BF",X"BF",X"BF",X"BF",X"C8",X"F3",X"C9",X"F3",
		X"CC",X"BF",X"BF",X"BF",X"BF",X"BF",X"AC",X"F3",X"AD",X"F3",X"BE",X"BF",X"BF",X"BF",X"BF",X"BF",
		X"8C",X"F3",X"8D",X"F3",X"CC",X"BF",X"BF",X"BF",X"A8",X"F3",X"A9",X"F3",X"BF",X"BF",X"BE",X"BF",
		X"BF",X"BF",X"88",X"F3",X"89",X"F3",X"BB",X"F3",X"CC",X"BF",X"BF",X"BF",X"ED",X"F3",X"BF",X"BF",
		X"BF",X"BF",X"BE",X"BF",X"BF",X"BF",X"CD",X"F3",X"BB",X"F3",X"BB",X"F3",X"CC",X"BF",X"5D",X"FA",
		X"E6",X"01",X"4C",X"A4",X"8F",X"3E",X"68",X"5F",X"CD",X"35",X"8F",X"35",X"00",X"1D",X"1C",X"01",
		X"10",X"0A",X"F2",X"86",X"A8",X"F3",X"E8",X"AC",X"41",X"F3",X"7A",X"AC",X"E6",X"F3",X"C2",X"AC",
		X"10",X"62",X"00",X"FB",X"F2",X"5C",X"9E",X"9B",X"53",X"45",X"8F",X"36",X"DC",X"4D",X"E0",X"4B",
		X"AE",X"83",X"DB",X"C1",X"A7",X"AE",X"8B",X"E0",X"60",X"40",X"AE",X"AB",X"8B",X"F0",X"8B",X"F1",
		X"DB",X"FB",X"BF",X"D8",X"8F",X"9C",X"CA",X"9E",X"E0",X"8B",X"E9",X"C8",X"F9",X"8B",X"5D",X"55",
		X"F8",X"8B",X"F9",X"8B",X"E0",X"08",X"9E",X"6A",X"C1",X"08",X"15",X"1D",X"B7",X"48",X"0D",X"8B",
		X"8B",X"8B",X"8B",X"B6",X"3C",X"0D",X"A2",X"52",X"F8",X"A3",X"3D",X"B5",X"4B",X"38",X"81",X"CE",
		X"A2",X"BD",X"D8",X"E6",X"69",X"9B",X"A3",X"BD",X"D8",X"A2",X"76",X"FC",X"4B",X"AE",X"9B",X"5C",
		X"0A",X"C2",X"53",X"A3",X"C6",X"D8",X"A3",X"E6",X"D8",X"C6",X"A3",X"DE",X"FC",X"5C",X"BF",X"D6",
		X"A2",X"4A",X"F8",X"D8",X"60",X"3E",X"E2",X"DA",X"AE",X"9E",X"84",X"69",X"7F",X"60",X"7F",X"E2",
		X"B7",X"AF",X"9B",X"5C",X"A6",X"BA",X"A2",X"B7",X"FC",X"4B",X"AF",X"DA",X"5C",X"CE",X"DB",X"A2",
		X"2F",X"F8",X"4B",X"E2",X"DB",X"A3",X"FD",X"D8",X"7D",X"38",X"CE",X"A2",X"B7",X"FC",X"4B",X"AE",
		X"FB",X"A2",X"BD",X"D8",X"4B",X"AE",X"EC",X"A2",X"0F",X"F8",X"4B",X"AE",X"E9",X"D9",X"8F",X"BA",
		X"D8",X"4D",X"A2",X"2E",X"F8",X"F8",X"06",X"AF",X"D2",X"A2",X"0E",X"F8",X"8B",X"F8",X"17",X"18",
		X"C0",X"AE",X"BB",X"4C",X"FD",X"60",X"9B",X"A7",X"DA",X"8B",X"8B",X"8B",X"E0",X"69",X"DA",X"60",
		X"DF",X"AF",X"DF",X"E2",X"9F",X"A3",X"2F",X"F8",X"0D",X"8B",X"8B",X"8B",X"8B",X"FA",X"BF",X"A2",
		X"B7",X"FC",X"4B",X"AF",X"B7",X"A2",X"BD",X"D8",X"4B",X"AF",X"CF",X"4C",X"D0",X"69",X"C2",X"60",
		X"FF",X"A7",X"BB",X"FA",X"3F",X"E0",X"0E",X"C1",X"69",X"DA",X"E6",X"FA",X"BF",X"18",X"E0",X"AE",
		X"FF",X"FA",X"3F",X"71",X"BB",X"4B",X"38",X"8C",X"CE",X"60",X"FB",X"38",X"E8",X"CE",X"07",X"C1",
		X"8B",X"B7",X"72",X"E2",X"9F",X"A3",X"C6",X"D8",X"A3",X"E6",X"D8",X"5C",X"BF",X"D6",X"A2",X"2F",
		X"F8",X"4B",X"E2",X"FB",X"A3",X"FD",X"D8",X"7D",X"38",X"CE",X"A2",X"C2",X"D8",X"4B",X"AE",X"9E",
		X"18",X"C1",X"AF",X"DF",X"E2",X"F3",X"5C",X"A6",X"BA",X"E2",X"BB",X"A3",X"C6",X"D8",X"A3",X"E6",
		X"D8",X"5C",X"BF",X"D6",X"A2",X"C2",X"D8",X"4B",X"AE",X"9E",X"18",X"C1",X"AF",X"DF",X"E2",X"93",
		X"5C",X"A6",X"BA",X"05",X"68",X"9F",X"45",X"D0",X"DB",X"1B",X"79",X"9B",X"D1",X"F2",X"9B",X"FB",
		X"9B",X"5D",X"55",X"80",X"A3",X"C6",X"D8",X"A0",X"A3",X"E6",X"D8",X"5C",X"BF",X"D6",X"A2",X"C2",
		X"D8",X"69",X"25",X"D8",X"60",X"2F",X"E2",X"97",X"AE",X"DB",X"84",X"60",X"37",X"E2",X"B3",X"AF",
		X"9B",X"5C",X"A6",X"BA",X"15",X"1D",X"F7",X"F6",X"B7",X"51",X"A2",X"2F",X"F8",X"4B",X"E2",X"DF",
		X"A3",X"FD",X"D8",X"7D",X"38",X"CE",X"A2",X"B7",X"FC",X"4B",X"AF",X"BE",X"E2",X"9E",X"A3",X"BF",
		X"FC",X"5C",X"DE",X"DF",X"FB",X"9E",X"5C",X"AA",X"EA",X"A3",X"3D",X"B5",X"B7",X"24",X"5C",X"8F",
		X"9B",X"05",X"19",X"16",X"8A",X"D4",X"C5",X"D2",X"49",X"41",X"CC",X"85",X"CC",X"68",X"37",X"CC",
		X"0B",X"58",X"6A",X"13",X"22",X"3B",X"7D",X"72",X"37",X"1E",X"36",X"A4",X"5F",X"22",X"B5",X"34",
		X"27",X"A9",X"94",X"1E",X"6C",X"E1",X"4A",X"41",X"8D",X"E2",X"9F",X"19",X"52",X"EE",X"E2",X"5F",
		X"19",X"52",X"EE",X"05",X"53",X"A3",X"C2",X"FC",X"E6",X"A3",X"2A",X"FC",X"8F",X"DB",X"DC",X"A2",
		X"FF",X"DC",X"60",X"9F",X"AE",X"9B",X"8F",X"BA",X"DC",X"F1",X"53",X"D8",X"4C",X"C8",X"D0",X"E0",
		X"D9",X"A1",X"80",X"5C",X"CA",X"DF",X"5C",X"8C",X"DB",X"A2",X"B7",X"FC",X"4B",X"AF",X"BE",X"E2",
		X"9E",X"A3",X"BF",X"FC",X"5C",X"DE",X"DF",X"5C",X"63",X"DB",X"E2",X"FF",X"5C",X"A6",X"BA",X"5C",
		X"A6",X"9B",X"53",X"A3",X"2F",X"F8",X"A2",X"FF",X"DC",X"8F",X"BD",X"FC",X"60",X"9F",X"AE",X"9B",
		X"8F",X"9D",X"FC",X"E3",X"9F",X"53",X"A3",X"2A",X"FC",X"1C",X"A2",X"72",X"F8",X"4B",X"3C",X"05",
		X"05",X"5C",X"63",X"DB",X"A2",X"FD",X"D8",X"5C",X"A6",X"BA",X"5C",X"B1",X"9B",X"53",X"A3",X"C2",
		X"FC",X"E6",X"A3",X"2A",X"FC",X"A3",X"2F",X"F8",X"A2",X"FF",X"DC",X"8F",X"BD",X"FC",X"97",X"0D",
		X"DC",X"9F",X"CC",X"F8",X"60",X"9F",X"AE",X"9E",X"8F",X"9D",X"FC",X"97",X"CB",X"F8",X"9F",X"E5",
		X"F8",X"E3",X"BF",X"5D",X"8F",X"B7",X"DC",X"FB",X"F9",X"E0",X"B3",X"8B",X"93",X"B7",X"20",X"15",
		X"A2",X"2B",X"F8",X"B3",X"93",X"8F",X"35",X"F8",X"FB",X"FB",X"E0",X"B3",X"5D",X"9F",X"9A",X"BF",
		X"9E",X"1D",X"93",X"B7",X"45",X"53",X"A3",X"2A",X"FC",X"1C",X"A2",X"C4",X"F8",X"4B",X"3C",X"8F",
		X"FA",X"FC",X"C7",X"3D",X"A2",X"C4",X"F8",X"C1",X"5C",X"8F",X"9B",X"1C",X"A2",X"E6",X"D8",X"60",
		X"BB",X"AE",X"88",X"60",X"9F",X"AE",X"90",X"4D",X"E0",X"60",X"37",X"AF",X"9E",X"4D",X"8B",X"8B",
		X"E8",X"EB",X"DC",X"18",X"62",X"0D",X"97",X"20",X"40",X"96",X"F9",X"A2",X"0E",X"F8",X"26",X"FB",
		X"BF",X"A6",X"9F",X"FF",X"8B",X"8B",X"8B",X"E3",X"E4",X"E2",X"9B",X"18",X"BD",X"AE",X"BB",X"4C",
		X"FD",X"D8",X"A2",X"E6",X"D8",X"71",X"9B",X"D0",X"DB",X"DB",X"1B",X"F3",X"BF",X"D0",X"8F",X"BC",
		X"D8",X"96",X"08",X"E2",X"E4",X"B3",X"93",X"E2",X"FA",X"B3",X"93",X"84",X"B3",X"93",X"53",X"B3",
		X"93",X"B3",X"93",X"0D",X"8A",X"A1",X"8A",X"81",X"8F",X"72",X"F8",X"C7",X"8F",X"A5",X"D8",X"E7",
		X"A4",X"1C",X"8B",X"A2",X"3B",X"F8",X"C1",X"FB",X"FE",X"97",X"E9",X"D8",X"B6",X"FA",X"8B",X"E3",
		X"F7",X"A2",X"0B",X"F8",X"DB",X"DB",X"79",X"B6",X"D9",X"97",X"88",X"D8",X"8A",X"8A",X"A4",X"B3",
		X"93",X"53",X"B3",X"93",X"B3",X"93",X"B3",X"93",X"E2",X"FE",X"B3",X"93",X"A1",X"8A",X"81",X"8A",
		X"A5",X"1C",X"4D",X"A2",X"E6",X"D8",X"60",X"BB",X"AE",X"DC",X"60",X"9F",X"AE",X"E3",X"8A",X"F1",
		X"8A",X"F0",X"92",X"92",X"92",X"92",X"B2",X"71",X"BB",X"B3",X"92",X"81",X"8B",X"A1",X"8A",X"8A",
		X"8A",X"8A",X"69",X"3F",X"AE",X"F6",X"E0",X"60",X"AF",X"A7",X"D3",X"53",X"8B",X"8B",X"C1",X"8B",
		X"8B",X"8B",X"C1",X"8F",X"52",X"F8",X"C7",X"8F",X"A5",X"D8",X"C7",X"AF",X"DF",X"E2",X"B6",X"5C",
		X"A6",X"BA",X"0D",X"1C",X"5C",X"86",X"CA",X"AF",X"04",X"E3",X"BA",X"8A",X"E3",X"3F",X"8A",X"97",
		X"B5",X"8B",X"A1",X"8A",X"81",X"B6",X"08",X"5C",X"86",X"CA",X"AF",X"69",X"A2",X"7F",X"F8",X"C1",
		X"8A",X"53",X"C1",X"8A",X"8A",X"8A",X"C1",X"B6",X"14",X"8A",X"F1",X"8A",X"F0",X"92",X"92",X"92",
		X"92",X"92",X"81",X"8B",X"A1",X"8B",X"8B",X"C7",X"1C",X"D4",X"CA",X"ED",X"CA",X"88",X"CA",X"A4",
		X"CA",X"3E",X"CA",X"0F",X"CA",X"2E",X"CA",X"ED",X"CA",X"26",X"CA",X"66",X"CA",X"BB",X"60",X"40",
		X"FB",X"70",X"40",X"FB",X"BB",X"40",X"40",X"FF",X"50",X"40",X"FF",X"FF",X"BF",X"BF",X"FF",X"2D",
		X"40",X"FF",X"40",X"40",X"FF",X"50",X"40",X"FF",X"DF",X"44",X"40",X"FE",X"46",X"40",X"FE",X"60",
		X"40",X"FA",X"62",X"40",X"BA",X"2D",X"40",X"7B",X"BE",X"44",X"40",X"FF",X"54",X"40",X"FF",X"60",
		X"40",X"FF",X"70",X"40",X"FF",X"44",X"9B",X"D3",X"54",X"9B",X"D3",X"60",X"9B",X"D3",X"70",X"9B",
		X"D3",X"BB",X"60",X"40",X"FE",X"70",X"40",X"FE",X"DF",X"60",X"40",X"B2",X"70",X"40",X"B2",X"40",
		X"40",X"F2",X"50",X"40",X"F2",X"BF",X"BF",X"B2",X"9F",X"44",X"40",X"9A",X"9F",X"44",X"40",X"9A",
		X"01",X"8F",X"D4",X"CA",X"97",X"F3",X"D9",X"9F",X"B7",X"C2",X"19",X"4B",X"E3",X"C6",X"A7",X"E0",
		X"A7",X"1D",X"A7",X"BE",X"87",X"D8",X"87",X"32",X"87",X"28",X"87",X"83",X"A3",X"1F",X"A3",X"78",
		X"A3",X"F2",X"83",X"E8",X"83",X"3D",X"83",X"97",X"E7",X"89",X"E7",X"07",X"E7",X"BB",X"C7",X"D8",
		X"C7",X"52",X"C7",X"00",X"CA",X"98",X"1A",X"0D",X"19",X"0F",X"96",X"17",X"3B",X"7A",X"5B",X"07",
		X"D7",X"5C",X"31",X"16",X"13",X"56",X"77",X"33",X"7A",X"7B",X"50",X"12",X"32",X"1F",X"53",X"73",
		X"27",X"32",X"59",X"9B",X"17",X"72",X"35",X"3E",X"5F",X"18",X"12",X"32",X"32",X"5A",X"17",X"31",
		X"FF",X"32",X"52",X"1F",X"72",X"35",X"7E",X"7B",X"18",X"12",X"32",X"36",X"77",X"37",X"1B",X"36",
		X"1C",X"7E",X"1F",X"7A",X"32",X"77",X"DF",X"23",X"BF",X"BB",X"16",X"7B",X"7A",X"13",X"5F",X"18",
		X"56",X"73",X"36",X"1F",X"B7",X"93",X"03",X"7F",X"1C",X"7E",X"7F",X"18",X"3A",X"3D",X"B6",X"32",
		X"3D",X"5A",X"32",X"51",X"FB",X"72",X"35",X"7E",X"7B",X"18",X"3A",X"32",X"36",X"1B",X"35",X"BB",
		X"03",X"32",X"1C",X"7E",X"7B",X"18",X"12",X"16",X"77",X"32",X"36",X"32",X"92",X"F7",X"33",X"74",
		X"7E",X"5F",X"18",X"3A",X"32",X"3F",X"13",X"2F",X"77",X"B3",X"11",X"32",X"1C",X"7E",X"33",X"5F",
		X"18",X"3A",X"17",X"27",X"57",X"3D",X"97",X"73",X"52",X"1F",X"72",X"35",X"7E",X"7F",X"18",X"12",
		X"B3",X"16",X"32",X"1F",X"DB",X"5A",X"43",X"3B",X"72",X"35",X"7E",X"1F",X"7A",X"D3",X"76",X"5A",
		X"BF",X"27",X"32",X"15",X"1B",X"7A",X"5F",X"50",X"56",X"77",X"31",X"73",X"32",X"16",X"DB",X"5A",
		X"03",X"57",X"1C",X"3E",X"7F",X"18",X"12",X"B2",X"7F",X"17",X"33",X"27",X"32",X"03",X"DF",X"74",
		X"7E",X"17",X"7F",X"7A",X"7F",X"16",X"5F",X"5A",X"30",X"3B",X"5A",X"FB",X"57",X"1B",X"7A",X"5F",
		X"50",X"3A",X"32",X"3F",X"DB",X"7C",X"73",X"72",X"35",X"3A",X"11",X"32",X"74",X"3E",X"7B",X"18",
		X"3A",X"96",X"75",X"1F",X"32",X"07",X"77",X"57",X"03",X"97",X"1C",X"7E",X"7F",X"18",X"56",X"B2",
		X"5B",X"D3",X"5C",X"B6",X"3F",X"32",X"9B",X"77",X"33",X"1C",X"7E",X"1F",X"7A",X"32",X"1F",X"17",
		X"5A",X"30",X"BB",X"5A",X"33",X"15",X"32",X"7A",X"13",X"7F",X"18",X"56",X"BF",X"DB",X"57",X"3D",
		X"5A",X"1F",X"43",X"B6",X"72",X"35",X"7E",X"7B",X"18",X"3A",X"32",X"3F",X"7B",X"11",X"5A",X"77",
		X"1B",X"12",X"F7",X"1C",X"7E",X"7F",X"18",X"12",X"3D",X"BB",X"17",X"1D",X"5A",X"7F",X"33",X"03",
		X"32",X"1C",X"7E",X"7B",X"18",X"3A",X"32",X"77",X"DF",X"75",X"5A",X"3F",X"11",X"DF",X"1C",X"7E",
		X"7F",X"18",X"12",X"75",X"73",X"53",X"1D",X"5A",X"17",X"77",X"83",X"77",X"32",X"1C",X"7E",X"33",
		X"7F",X"18",X"12",X"F7",X"5B",X"57",X"23",X"DA",X"53",X"43",X"5B",X"72",X"35",X"7E",X"5F",X"7A",
		X"DA",X"32",X"3B",X"5C",X"1F",X"A3",X"5A",X"32",X"5C",X"55",X"32",X"5A",X"7A",X"7B",X"50",X"12",
		X"16",X"32",X"F3",X"32",X"23",X"5A",X"B6",X"5B",X"17",X"72",X"35",X"3E",X"1F",X"7A",X"32",X"3B",
		X"5C",X"3F",X"A3",X"5A",X"32",X"5C",X"15",X"B2",X"7A",X"5F",X"50",X"12",X"7B",X"23",X"7B",X"B2",
		X"2B",X"5A",X"77",X"77",X"DB",X"13",X"33",X"72",X"35",X"3E",X"17",X"7F",X"18",X"56",X"F7",X"DB",
		X"5A",X"B2",X"3F",X"5A",X"73",X"11",X"D7",X"74",X"7E",X"7B",X"18",X"12",X"32",X"3B",X"53",X"5A",
		X"47",X"5A",X"1B",X"93",X"5B",X"1C",X"3A",X"1E",X"7E",X"7B",X"18",X"3A",X"17",X"15",X"32",X"5A",
		X"1D",X"5A",X"7F",X"36",X"4A",X"FF",X"72",X"35",X"3A",X"1E",X"7E",X"7B",X"18",X"12",X"32",X"32",
		X"3B",X"5A",X"2F",X"5A",X"93",X"49",X"77",X"33",X"1C",X"3A",X"1E",X"7E",X"7B",X"18",X"3A",X"1F",
		X"75",X"32",X"5A",X"B6",X"5F",X"5A",X"93",X"FB",X"74",X"7E",X"13",X"5F",X"18",X"56",X"5B",X"16",
		X"5A",X"93",X"57",X"77",X"33",X"52",X"17",X"72",X"35",X"7E",X"5F",X"7A",X"5A",X"32",X"7F",X"1C",
		X"56",X"F7",X"5A",X"36",X"47",X"3B",X"B3",X"7A",X"7F",X"7A",X"53",X"F6",X"FF",X"5A",X"32",X"22",
		X"1C",X"56",X"5A",X"55",X"DF",X"53",X"7A",X"7F",X"7A",X"D7",X"0F",X"73",X"73",X"77",X"34",X"5A",
		X"32",X"9D",X"1C",X"56",X"5A",X"7A",X"7F",X"50",X"12",X"F7",X"7B",X"BF",X"15",X"1B",X"5A",X"11",
		X"32",X"74",X"3E",X"33",X"7B",X"18",X"56",X"16",X"3F",X"BF",X"31",X"5A",X"F3",X"5B",X"36",X"72",
		X"35",X"7E",X"7B",X"18",X"3A",X"BB",X"BB",X"32",X"5C",X"5A",X"BB",X"32",X"5A",X"5C",X"9B",X"32",
		X"53",X"1C",X"7E",X"7F",X"7A",X"32",X"74",X"1B",X"5C",X"32",X"14",X"5A",X"32",X"5C",X"14",X"5B",
		X"32",X"7A",X"7B",X"50",X"3A",X"9F",X"BB",X"32",X"5C",X"5A",X"BB",X"32",X"5A",X"5C",X"9B",X"32",
		X"FF",X"1C",X"3E",X"5F",X"18",X"12",X"7B",X"77",X"32",X"34",X"5A",X"32",X"83",X"77",X"93",X"74",
		X"7E",X"17",X"7F",X"18",X"56",X"B3",X"93",X"5A",X"39",X"5C",X"5A",X"D7",X"43",X"17",X"72",X"35",
		X"7E",X"7F",X"7A",X"32",X"74",X"5C",X"5B",X"32",X"14",X"5C",X"32",X"5B",X"14",X"5C",X"32",X"7A",
		X"5F",X"50",X"12",X"9B",X"07",X"32",X"5A",X"39",X"1F",X"5C",X"32",X"03",X"F3",X"74",X"3E",X"7F",
		X"7A",X"5A",X"9F",X"7F",X"DF",X"5C",X"31",X"32",X"5B",X"14",X"5C",X"32",X"7A",X"5F",X"50",X"56",
		X"3B",X"0B",X"5A",X"5A",X"77",X"5A",X"30",X"5A",X"33",X"32",X"12",X"FB",X"1C",X"3E",X"13",X"7B",
		X"18",X"12",X"16",X"32",X"9B",X"1F",X"3D",X"5A",X"D3",X"4B",X"73",X"33",X"72",X"35",X"7E",X"3B",
		X"7A",X"5A",X"A9",X"1C",X"56",X"5B",X"5A",X"DB",X"BB",X"32",X"5B",X"5A",X"8F",X"DB",X"5C",X"5A",
		X"7A",X"7F",X"7A",X"32",X"36",X"32",X"75",X"5C",X"32",X"16",X"32",X"7A",X"7B",X"50",X"12",X"32",
		X"2F",X"5C",X"32",X"BC",X"F7",X"5A",X"77",X"32",X"83",X"5C",X"32",X"74",X"3E",X"7F",X"7A",X"32",
		X"30",X"5A",X"77",X"5F",X"84",X"72",X"35",X"56",X"FB",X"36",X"14",X"5A",X"32",X"7A",X"33",X"5F",
		X"18",X"12",X"5A",X"74",X"5A",X"5A",X"93",X"2B",X"77",X"B3",X"5A",X"C3",X"5A",X"5A",X"72",X"35",
		X"7E",X"7B",X"18",X"12",X"B2",X"32",X"5C",X"5A",X"9F",X"13",X"5A",X"5C",X"51",X"32",X"72",X"35",
		X"7E",X"5B",X"18",X"56",X"77",X"32",X"76",X"5C",X"B2",X"14",X"5C",X"32",X"5C",X"01",X"77",X"B2",
		X"74",X"7E",X"7B",X"18",X"12",X"32",X"36",X"57",X"96",X"F3",X"32",X"5C",X"51",X"32",X"72",X"35",
		X"7E",X"5F",X"18",X"56",X"5F",X"32",X"36",X"7B",X"77",X"1B",X"03",X"32",X"74",X"7E",X"17",X"1F",
		X"7A",X"5A",X"11",X"13",X"77",X"33",X"65",X"1C",X"56",X"1F",X"56",X"5A",X"BB",X"7A",X"7B",X"50",
		X"12",X"32",X"46",X"77",X"5C",X"BF",X"5F",X"23",X"32",X"5C",X"83",X"5A",X"32",X"74",X"3E",X"7B",
		X"18",X"3A",X"53",X"F7",X"32",X"D7",X"C7",X"5C",X"1B",X"5A",X"32",X"1B",X"FF",X"1C",X"7E",X"7B",
		X"18",X"12",X"32",X"2B",X"3F",X"5C",X"17",X"AF",X"73",X"5A",X"32",X"D0",X"1C",X"56",X"DB",X"72",
		X"35",X"7E",X"7F",X"7A",X"7B",X"BB",X"32",X"5C",X"BB",X"31",X"32",X"36",X"87",X"5C",X"32",X"7A",
		X"13",X"5F",X"18",X"56",X"7B",X"32",X"DA",X"5B",X"1D",X"5A",X"96",X"5A",X"11",X"13",X"74",X"7E",
		X"5F",X"18",X"3A",X"5A",X"23",X"32",X"5C",X"BB",X"32",X"5C",X"32",X"0B",X"77",X"33",X"1C",X"7E",
		X"7B",X"18",X"12",X"32",X"56",X"5C",X"96",X"5A",X"55",X"32",X"5C",X"32",X"52",X"5A",X"77",X"1C",
		X"7E",X"5F",X"18",X"3A",X"32",X"56",X"DF",X"5C",X"32",X"76",X"5C",X"D3",X"83",X"1B",X"32",X"74",
		X"7E",X"7B",X"18",X"12",X"53",X"34",X"7F",X"17",X"F7",X"32",X"57",X"59",X"73",X"97",X"72",X"35",
		X"7E",X"33",X"7B",X"18",X"3A",X"17",X"F6",X"17",X"FF",X"5C",X"14",X"D3",X"5C",X"DF",X"10",X"5C",
		X"DB",X"1C",X"7E",X"7B",X"18",X"3A",X"16",X"BB",X"32",X"5C",X"32",X"2F",X"5C",X"32",X"83",X"5C",
		X"32",X"74",X"7E",X"5B",X"18",X"56",X"77",X"32",X"76",X"5C",X"32",X"14",X"5C",X"32",X"5C",X"51",
		X"32",X"72",X"35",X"7E",X"7B",X"18",X"12",X"32",X"2F",X"5C",X"32",X"A3",X"5C",X"32",X"5C",X"9B",
		X"32",X"F3",X"1C",X"7E",X"7F",X"7A",X"32",X"14",X"5A",X"32",X"5A",X"55",X"32",X"5A",X"32",X"56",
		X"5A",X"B6",X"7A",X"17",X"7F",X"18",X"56",X"B2",X"5A",X"5A",X"5A",X"1D",X"DA",X"5A",X"5A",X"03",
		X"5A",X"74",X"7E",X"7B",X"18",X"12",X"32",X"47",X"5C",X"53",X"1B",X"5D",X"D3",X"1C",X"56",X"B6",
		X"03",X"32",X"74",X"7E",X"7F",X"7A",X"32",X"14",X"5C",X"32",X"5C",X"75",X"32",X"32",X"54",X"5C",
		X"5A",X"5A",X"7A",X"7B",X"50",X"12",X"32",X"2F",X"5C",X"32",X"31",X"93",X"33",X"83",X"5C",X"32",
		X"74",X"3E",X"5F",X"18",X"12",X"32",X"76",X"5C",X"DF",X"BF",X"3F",X"32",X"83",X"5C",X"B2",X"74",
		X"7E",X"13",X"5F",X"7A",X"BF",X"5A",X"28",X"72",X"35",X"3A",X"16",X"57",X"55",X"17",X"5A",X"5A",
		X"16",X"93",X"7A",X"7B",X"50",X"12",X"32",X"67",X"5A",X"5B",X"A3",X"5C",X"32",X"5C",X"D3",X"32",
		X"77",X"1C",X"3E",X"7B",X"18",X"12",X"32",X"2F",X"5C",X"32",X"A3",X"5C",X"32",X"D7",X"19",X"5C",
		X"B6",X"1C",X"7E",X"7B",X"18",X"12",X"32",X"2F",X"5C",X"32",X"B2",X"7F",X"9F",X"3B",X"03",X"32",
		X"74",X"7E",X"7B",X"18",X"12",X"32",X"66",X"1C",X"56",X"DF",X"96",X"53",X"5F",X"1B",X"03",X"32",
		X"74",X"7E",X"33",X"7B",X"18",X"3A",X"BF",X"A3",X"5B",X"5C",X"36",X"BF",X"B6",X"5C",X"59",X"73",
		X"53",X"72",X"35",X"7E",X"1F",X"7A",X"32",X"16",X"32",X"5C",X"75",X"32",X"32",X"55",X"5C",X"BF",
		X"7A",X"7B",X"50",X"3A",X"5A",X"AB",X"5A",X"5A",X"5A",X"5A",X"AB",X"5A",X"DA",X"5A",X"5A",X"83",
		X"5A",X"32",X"74",X"3E",X"7F",X"7A",X"32",X"34",X"5C",X"1F",X"87",X"F7",X"13",X"7F",X"0F",X"77",
		X"33",X"7A",X"3B",X"7A",X"3B",X"14",X"5C",X"32",X"9B",X"32",X"7B",X"7B",X"16",X"5F",X"7A",X"17",
		X"7F",X"18",X"3A",X"E7",X"73",X"D3",X"17",X"2B",X"7F",X"5C",X"5A",X"8B",X"DA",X"5A",X"5A",X"1C",
		X"7E",X"7F",X"7A",X"32",X"15",X"5C",X"32",X"76",X"5C",X"32",X"14",X"5C",X"32",X"7A",X"7F",X"7A",
		X"D7",X"A3",X"5C",X"32",X"5C",X"BB",X"32",X"5C",X"32",X"47",X"D7",X"17",X"7A",X"5F",X"7A",X"9F",
		X"72",X"A1",X"35",X"3A",X"32",X"5C",X"D5",X"77",X"32",X"33",X"5C",X"55",X"16",X"36",X"7A",X"7B",
		X"50",X"3A",X"7B",X"23",X"32",X"5C",X"BB",X"32",X"5A",X"B6",X"83",X"5A",X"32",X"74",X"3E",X"13",
		X"5F",X"7A",X"5A",X"BF",X"10",X"5C",X"D3",X"73",X"72",X"A9",X"35",X"3A",X"DB",X"5C",X"3B",X"55",
		X"7F",X"5A",X"7A",X"7B",X"50",X"3A",X"16",X"03",X"32",X"1C",X"56",X"D1",X"77",X"32",X"77",X"72",
		X"35",X"81",X"56",X"77",X"32",X"74",X"3E",X"5F",X"18",X"56",X"32",X"76",X"5C",X"57",X"A3",X"97",
		X"32",X"5C",X"9B",X"32",X"33",X"1C",X"7E",X"7B",X"18",X"12",X"32",X"2F",X"5C",X"32",X"AF",X"5C",
		X"77",X"93",X"83",X"33",X"32",X"74",X"7E",X"5F",X"7A",X"5A",X"32",X"16",X"32",X"5C",X"75",X"32",
		X"7B",X"54",X"BF",X"5F",X"5A",X"7A",X"3B",X"1F",X"D2",X"E3",X"CB",X"E3",X"CA",X"E3",X"C3",X"E3",
		X"C2",X"E3",X"D9",X"E3",X"D8",X"E3",X"D1",X"E3",X"D0",X"E3",X"C9",X"E3",X"C8",X"E3",X"C1",X"E3",
		X"C0",X"E3",X"5B",X"E3",X"5A",X"E3",X"53",X"E3",X"52",X"E3",X"10",X"F3",X"19",X"2B",X"9F",X"FF",
		X"F3",X"DA",X"25",X"BD",X"B7",X"BE",X"FF",X"DF",X"D7",X"FA",X"2D",X"E6",X"AF",X"BA",X"FF",X"FB",
		X"F7",X"DE",X"35",X"A6",X"A7",X"FE",X"FF",X"DB",X"93",X"FE",X"3D",X"E7",X"BD",X"FA",X"FF",X"BE",
		X"B3",X"9A",X"27",X"A7",X"B5",X"B7",X"FF",X"9E",X"97",X"BA",X"2F",X"EE",X"AD",X"F7",X"DF",X"BA",
		X"B7",X"9E",X"37",X"AE",X"A5",X"B6",X"DF",X"9A",X"DA",X"BE",X"3F",X"EB",X"3F",X"F6",X"DF",X"DE",
		X"FA",X"DB",X"A5",X"EF",X"37",X"AF",X"DF",X"DA",X"DE",X"FB",X"AD",X"AB",X"2F",X"EF",X"DF",X"B3",
		X"FE",X"FB",X"B5",X"AF",X"27",X"AE",X"FB",X"F3",X"9A",X"FB",X"BD",X"F2",X"3D",X"EE",X"FB",X"F2",
		X"BA",X"DF",X"A7",X"F6",X"35",X"A7",X"FB",X"CE",X"9E",X"DF",X"AF",X"B2",X"2D",X"E7",X"FB",X"B0",
		X"BE",X"DF",X"B7",X"B6",X"25",X"A6",X"DB",X"9B",X"3F",X"9F",X"D8",X"96",X"E7",X"BA",X"FF",X"DF",
		X"3F",X"9F",X"BC",X"B6",X"EE",X"DF",X"FF",X"55",X"08",X"8F",X"BF",X"BF",X"B2",X"55",X"F3",X"BF",
		X"D0",X"96",X"15",X"92",X"B7",X"61",X"E2",X"FB",X"A3",X"3D",X"B5",X"A3",X"BA",X"FC",X"E6",X"E6",
		X"A3",X"9A",X"FC",X"DE",X"AF",X"69",X"15",X"96",X"E4",X"69",X"C2",X"C9",X"0C",X"A2",X"82",X"FC",
		X"60",X"9F",X"AE",X"EB",X"54",X"8F",X"32",X"FC",X"8F",X"2B",X"FC",X"97",X"B8",X"FC",X"FB",X"9B",
		X"E0",X"B3",X"8A",X"92",X"B7",X"20",X"5C",X"6E",X"86",X"A2",X"53",X"FC",X"4B",X"AF",X"BE",X"5C",
		X"CF",X"C3",X"5C",X"EE",X"C3",X"B6",X"FB",X"5C",X"EE",X"C3",X"5C",X"CF",X"C3",X"A2",X"32",X"FC",
		X"60",X"9F",X"3D",X"53",X"A3",X"32",X"FC",X"5C",X"37",X"A2",X"FB",X"67",X"5C",X"9E",X"9B",X"1C",
		X"A2",X"BA",X"FC",X"D9",X"97",X"98",X"FC",X"E0",X"B3",X"8B",X"93",X"B7",X"20",X"5C",X"A2",X"C3",
		X"53",X"5C",X"FC",X"BB",X"1C",X"8F",X"56",X"FC",X"E2",X"9F",X"B6",X"DF",X"8F",X"2F",X"FC",X"E2",
		X"BB",X"A3",X"37",X"FC",X"5C",X"25",X"9F",X"19",X"31",X"FF",X"A2",X"16",X"FC",X"60",X"BA",X"AE",
		X"FF",X"E6",X"A3",X"16",X"FC",X"54",X"8F",X"7F",X"FC",X"8F",X"98",X"FC",X"97",X"BC",X"FC",X"FB",
		X"9B",X"E0",X"B3",X"8B",X"93",X"B7",X"20",X"5C",X"6E",X"86",X"A2",X"53",X"FC",X"4B",X"3C",X"01",
		X"10",X"CD",X"F2",X"03",X"C7",X"89",X"F2",X"23",X"C7",X"75",X"F3",X"70",X"AC",X"D5",X"48",X"AC",
		X"29",X"F9",X"89",X"DA",X"A2",X"F1",X"D0",X"F5",X"32",X"41",X"F1",X"D0",X"F1",X"D0",X"F1",X"10",
		X"F3",X"00",X"5C",X"1E",X"C3",X"5C",X"91",X"86",X"1C",X"53",X"5C",X"FC",X"BB",X"E2",X"9E",X"5C",
		X"A6",X"BA",X"FB",X"E6",X"5C",X"9E",X"9B",X"5C",X"CE",X"FB",X"A3",X"33",X"FC",X"97",X"21",X"86",
		X"8F",X"7B",X"B9",X"5C",X"9C",X"FF",X"A2",X"37",X"FC",X"60",X"9F",X"E2",X"A3",X"AF",X"9F",X"C6",
		X"A3",X"5B",X"9D",X"E2",X"9E",X"5C",X"A6",X"9B",X"97",X"CF",X"A2",X"8F",X"2A",X"99",X"5C",X"9C",
		X"FF",X"97",X"CD",X"A2",X"8F",X"88",X"B9",X"5C",X"9C",X"FF",X"97",X"F6",X"A2",X"8F",X"B1",X"B9",
		X"5C",X"9C",X"FF",X"97",X"DE",X"A2",X"8F",X"30",X"B9",X"5C",X"9C",X"FF",X"E2",X"A7",X"A3",X"17",
		X"FC",X"5C",X"83",X"86",X"E2",X"F7",X"A3",X"13",X"FC",X"97",X"73",X"FC",X"E2",X"9F",X"A3",X"57",
		X"FC",X"E2",X"9D",X"B3",X"5C",X"DE",X"86",X"FB",X"E6",X"A3",X"BE",X"FC",X"5C",X"4D",X"A6",X"A2",
		X"33",X"FC",X"60",X"9F",X"3C",X"5C",X"F7",X"BB",X"18",X"C1",X"AF",X"82",X"A2",X"57",X"FC",X"69",
		X"9F",X"E2",X"BA",X"AE",X"BB",X"E2",X"D3",X"5C",X"A6",X"BA",X"A2",X"57",X"FC",X"8F",X"1E",X"FC",
		X"5F",X"C8",X"E4",X"78",X"BF",X"C9",X"B2",X"C1",X"A2",X"57",X"FC",X"60",X"9B",X"3C",X"E6",X"A3",
		X"57",X"FC",X"5C",X"F7",X"BB",X"18",X"C1",X"AF",X"9A",X"5C",X"4D",X"A6",X"A2",X"33",X"FC",X"60",
		X"9F",X"3C",X"B6",X"68",X"5C",X"DE",X"86",X"5C",X"F7",X"BB",X"18",X"D0",X"AF",X"9A",X"B2",X"C6",
		X"60",X"82",X"AF",X"BB",X"E2",X"B0",X"B3",X"B6",X"DA",X"5C",X"F7",X"BB",X"18",X"D9",X"AF",X"76",
		X"B2",X"E6",X"60",X"90",X"AF",X"BB",X"E2",X"E6",X"B3",X"5C",X"DE",X"86",X"A2",X"13",X"FC",X"60",
		X"FB",X"A6",X"DF",X"C6",X"C6",X"A3",X"13",X"FC",X"A3",X"77",X"FC",X"5C",X"F7",X"BB",X"A3",X"3D",
		X"B5",X"18",X"D0",X"AE",X"FE",X"18",X"D9",X"AE",X"BE",X"E2",X"F7",X"A3",X"13",X"FC",X"19",X"64",
		X"C3",X"A2",X"BE",X"FC",X"4B",X"AF",X"20",X"E2",X"9F",X"A3",X"BE",X"FC",X"B7",X"93",X"FB",X"E6",
		X"A2",X"17",X"FC",X"71",X"9F",X"CB",X"A3",X"17",X"FC",X"5C",X"83",X"86",X"A2",X"17",X"FC",X"4B",
		X"3C",X"8F",X"77",X"FC",X"C7",X"AF",X"7D",X"A2",X"13",X"FC",X"60",X"FB",X"A6",X"DF",X"C6",X"C6",
		X"A3",X"13",X"FC",X"C1",X"5C",X"F7",X"BB",X"18",X"D0",X"AF",X"9A",X"B2",X"C6",X"60",X"82",X"AF",
		X"BB",X"E2",X"B0",X"B3",X"B6",X"BE",X"B2",X"E6",X"60",X"90",X"AF",X"BB",X"E2",X"E6",X"B3",X"5C",
		X"DE",X"86",X"19",X"80",X"A6",X"A2",X"BE",X"FC",X"A3",X"3D",X"B5",X"4B",X"AF",X"41",X"E2",X"9F",
		X"A3",X"BE",X"FC",X"B7",X"D3",X"FB",X"E6",X"A2",X"17",X"FC",X"71",X"9F",X"CB",X"A3",X"17",X"FC",
		X"5C",X"83",X"86",X"4B",X"AE",X"9F",X"1C",X"E2",X"9F",X"A3",X"33",X"FC",X"1C",X"45",X"5D",X"4D",
		X"8F",X"B1",X"B9",X"A2",X"57",X"FC",X"60",X"BB",X"AF",X"9B",X"8F",X"B3",X"B9",X"60",X"9B",X"AF",
		X"9B",X"8F",X"31",X"9D",X"E2",X"DE",X"A3",X"BF",X"FC",X"A2",X"73",X"FC",X"5C",X"78",X"9B",X"0D",
		X"1D",X"05",X"1C",X"8F",X"B0",X"9D",X"45",X"53",X"A3",X"FB",X"FC",X"A2",X"12",X"FC",X"E6",X"60",
		X"DA",X"A6",X"BB",X"E2",X"9F",X"A3",X"12",X"FC",X"A3",X"BF",X"FC",X"A2",X"17",X"FC",X"5C",X"4B",
		X"9B",X"05",X"1C",X"9F",X"BA",X"BA",X"54",X"8F",X"F8",X"FC",X"8F",X"91",X"FC",X"97",X"F5",X"FC",
		X"A3",X"3D",X"B5",X"5D",X"FB",X"FB",X"4D",X"8F",X"DD",X"FC",X"B2",X"C1",X"93",X"8B",X"B7",X"20",
		X"0D",X"92",X"5C",X"6E",X"86",X"A2",X"53",X"FC",X"60",X"9F",X"AF",X"D6",X"FB",X"FB",X"E0",X"B3",
		X"8A",X"92",X"B7",X"20",X"8B",X"93",X"FB",X"FB",X"55",X"97",X"DD",X"FC",X"B2",X"C1",X"93",X"8B",
		X"B7",X"20",X"15",X"8A",X"93",X"93",X"93",X"93",X"93",X"93",X"55",X"97",X"FB",X"BF",X"96",X"54",
		X"96",X"15",X"1D",X"B7",X"02",X"FB",X"BA",X"DE",X"39",X"F1",X"86",X"1C",X"45",X"55",X"4D",X"8F",
		X"FB",X"FC",X"53",X"C1",X"A3",X"53",X"FC",X"97",X"B8",X"FC",X"B2",X"54",X"73",X"DF",X"CB",X"45",
		X"4B",X"AE",X"9B",X"E2",X"9F",X"C1",X"05",X"92",X"B2",X"54",X"72",X"FF",X"CB",X"45",X"4B",X"AE",
		X"9B",X"E2",X"9F",X"C1",X"05",X"92",X"B2",X"54",X"72",X"9B",X"CB",X"45",X"4B",X"AE",X"9B",X"E2",
		X"9F",X"C1",X"05",X"A6",X"9E",X"E0",X"4B",X"AE",X"DF",X"E2",X"9F",X"A3",X"53",X"FC",X"0D",X"15",
		X"05",X"1C",X"8A",X"65",X"01",X"30",X"05",X"15",X"24",X"77",X"10",X"11",X"09",X"30",X"05",X"8A",
		X"AA",X"34",X"2D",X"15",X"1C",X"05",X"30",X"77",X"77",X"77",X"57",X"8A",X"8A",X"8A",X"41",X"24",
		X"1D",X"0D",X"05",X"77",X"2D",X"05",X"21",X"24",X"8A",X"4D",X"8A",X"8A",X"8A",X"5D",X"08",X"77",
		X"08",X"77",X"08",X"8A",X"8A",X"8A",X"5D",X"0D",X"09",X"20",X"05",X"77",X"39",X"09",X"1C",X"10",
		X"24",X"1D",X"11",X"19",X"77",X"8A",X"71",X"04",X"34",X"77",X"8A",X"5D",X"09",X"30",X"77",X"8A",
		X"7D",X"25",X"09",X"00",X"29",X"8A",X"5D",X"8A",X"AA",X"24",X"09",X"77",X"10",X"05",X"2D",X"05",
		X"11",X"24",X"77",X"8A",X"AA",X"3D",X"1D",X"24",X"77",X"8A",X"65",X"34",X"04",X"29",X"11",X"3D",
		X"77",X"8A",X"5D",X"8A",X"8A",X"2D",X"05",X"24",X"24",X"05",X"30",X"10",X"6B",X"8A",X"AA",X"24",
		X"09",X"77",X"05",X"29",X"24",X"05",X"30",X"77",X"1D",X"29",X"1D",X"24",X"1D",X"15",X"2D",X"10",
		X"6B",X"8A",X"8A",X"8A",X"4D",X"05",X"3C",X"09",X"30",X"11",X"1D",X"10",X"24",X"10",X"8A",X"8A",
		X"53",X"5C",X"D5",X"BB",X"5C",X"CE",X"FB",X"97",X"1B",X"A2",X"8F",X"E9",X"B9",X"5C",X"9C",X"FF",
		X"9F",X"9F",X"BA",X"97",X"95",X"FC",X"8F",X"9E",X"99",X"4D",X"5C",X"39",X"A2",X"8F",X"FB",X"BF",
		X"96",X"08",X"0D",X"8B",X"8B",X"A2",X"16",X"FC",X"06",X"3C",X"84",X"79",X"9F",X"CB",X"D8",X"B7",
		X"2C",X"1C",X"5D",X"55",X"E2",X"9F",X"A3",X"FB",X"FC",X"E6",X"A3",X"BF",X"FC",X"84",X"5C",X"4B",
		X"9B",X"E2",X"EA",X"5C",X"78",X"9B",X"9F",X"3D",X"40",X"9E",X"E2",X"9F",X"A3",X"FB",X"FC",X"E2",
		X"9E",X"A3",X"BF",X"FC",X"5C",X"5E",X"9B",X"9F",X"AD",X"40",X"9E",X"E2",X"FF",X"A3",X"BF",X"FC",
		X"FB",X"9B",X"92",X"B2",X"5C",X"78",X"9B",X"5D",X"9F",X"BD",X"BF",X"9E",X"1D",X"B7",X"01",X"15",
		X"1D",X"1C",X"E2",X"9F",X"A3",X"B7",X"FC",X"A3",X"FF",X"DC",X"5C",X"61",X"9F",X"A2",X"3F",X"B5",
		X"18",X"C8",X"E2",X"9F",X"AE",X"9F",X"53",X"A3",X"97",X"FC",X"9F",X"F7",X"BF",X"F3",X"9F",X"E2",
		X"B7",X"5C",X"C6",X"82",X"9F",X"9F",X"9F",X"D1",X"E2",X"97",X"5C",X"C6",X"82",X"5C",X"37",X"A2",
		X"5C",X"38",X"FB",X"5C",X"1D",X"C6",X"FA",X"BE",X"5C",X"19",X"BB",X"B6",X"54",X"A3",X"BE",X"DC",
		X"A0",X"A3",X"76",X"FC",X"E2",X"9F",X"8F",X"FF",X"DC",X"C1",X"8B",X"A5",X"8B",X"85",X"A3",X"BD",
		X"FC",X"A3",X"B9",X"FC",X"5C",X"56",X"EF",X"01",X"10",X"B1",X"98",X"24",X"2A",X"C0",X"46",X"51",
		X"98",X"0F",X"98",X"D7",X"00",X"53",X"8F",X"93",X"FC",X"97",X"FF",X"BF",X"C1",X"96",X"B7",X"64",
		X"5C",X"00",X"DF",X"5C",X"38",X"FB",X"53",X"A3",X"4F",X"F8",X"E2",X"BA",X"A3",X"BF",X"FC",X"5C",
		X"F7",X"DF",X"5C",X"11",X"DF",X"A2",X"B3",X"FC",X"60",X"9F",X"AE",X"FB",X"5C",X"F6",X"DF",X"5C",
		X"70",X"DF",X"E2",X"9F",X"A3",X"4F",X"F8",X"5C",X"C0",X"8A",X"53",X"1C",X"45",X"5D",X"4D",X"A2",
		X"E6",X"D8",X"DB",X"DB",X"FB",X"BF",X"D8",X"8F",X"93",X"FC",X"9E",X"E0",X"4B",X"AF",X"9C",X"4D",
		X"A2",X"DF",X"DC",X"4B",X"8F",X"DB",X"E6",X"AE",X"9E",X"60",X"9F",X"8F",X"69",X"E6",X"AE",X"BB",
		X"B6",X"60",X"18",X"96",X"9E",X"F8",X"8B",X"F9",X"0D",X"4D",X"8B",X"8B",X"85",X"8B",X"A5",X"0D",
		X"4D",X"8B",X"8B",X"F8",X"8B",X"F9",X"0D",X"01",X"10",X"53",X"F8",X"80",X"10",X"3C",X"00",X"80",
		X"4B",X"AE",X"66",X"4D",X"E6",X"C1",X"9B",X"8B",X"01",X"10",X"53",X"F8",X"80",X"10",X"3C",X"00",
		X"80",X"C1",X"9B",X"8B",X"85",X"8B",X"A5",X"0D",X"C7",X"AE",X"55",X"8B",X"E0",X"A3",X"C3",X"FC",
		X"5C",X"0D",X"BB",X"0D",X"1D",X"05",X"1C",X"96",X"E6",X"A9",X"E6",X"88",X"E6",X"E4",X"E6",X"13",
		X"E6",X"27",X"E6",X"59",X"E6",X"31",X"E6",X"54",X"E6",X"CD",X"7D",X"ED",X"4D",X"F9",X"7D",X"CD",
		X"7C",X"F9",X"7D",X"F2",X"6D",X"DD",X"7D",X"CD",X"7C",X"F9",X"7D",X"F5",X"6D",X"D9",X"7D",X"CD",
		X"7C",X"F9",X"7D",X"CC",X"6D",X"DD",X"7D",X"CD",X"7C",X"F9",X"7D",X"FB",X"6D",X"E5",X"49",X"ED",
		X"4D",X"F8",X"7D",X"F9",X"4D",X"FC",X"7D",X"E8",X"4D",X"F8",X"7D",X"F5",X"4D",X"F8",X"7D",X"FC",
		X"7C",X"CD",X"7D",X"F4",X"4D",X"F8",X"49",X"D9",X"7D",X"E0",X"6D",X"C8",X"7C",X"D8",X"7D",X"F3",
		X"6D",X"FD",X"C1",X"69",X"C9",X"6D",X"F9",X"6D",X"F9",X"69",X"FD",X"F8",X"4D",X"C8",X"6D",X"F1",
		X"4D",X"CC",X"6D",X"F9",X"7D",X"D4",X"6D",X"F8",X"49",X"F3",X"4D",X"FD",X"C9",X"4D",X"CD",X"6D",
		X"C8",X"75",X"CD",X"7D",X"F3",X"6D",X"C8",X"75",X"CD",X"7D",X"F7",X"4D",X"DC",X"6D",X"D4",X"4D",
		X"CD",X"7F",X"FD",X"CD",X"7D",X"E9",X"6D",X"C8",X"4D",X"C8",X"75",X"CD",X"7D",X"D0",X"6D",X"F8",
		X"49",X"FC",X"6D",X"F9",X"7D",X"DB",X"4D",X"C4",X"6D",X"F8",X"69",X"F9",X"7D",X"F3",X"6D",X"FD",
		X"DC",X"6D",X"C8",X"75",X"CD",X"7D",X"F8",X"4D",X"C8",X"75",X"CD",X"7D",X"EF",X"4D",X"E0",X"6D",
		X"C5",X"4D",X"CF",X"6D",X"CD",X"5F",X"FD",X"DC",X"7D",X"F5",X"6D",X"F5",X"4D",X"C8",X"75",X"F3",
		X"4D",X"FD",X"E9",X"7D",X"F5",X"6D",X"F5",X"4D",X"CC",X"75",X"F3",X"7D",X"FD",X"D9",X"7D",X"F5",
		X"6D",X"F5",X"4D",X"F3",X"75",X"FD",X"24",X"E6",X"8E",X"C6",X"A3",X"C6",X"C2",X"C6",X"F5",X"C6",
		X"C8",X"C6",X"7B",X"C6",X"53",X"C6",X"27",X"C6",X"CD",X"7D",X"FF",X"4D",X"FC",X"7C",X"FC",X"7D",
		X"F5",X"4D",X"FC",X"7C",X"FC",X"7D",X"F5",X"4D",X"FC",X"7C",X"FC",X"7D",X"C5",X"4D",X"F8",X"49",
		X"F4",X"6D",X"F8",X"49",X"DC",X"6D",X"CD",X"7D",X"FC",X"7C",X"FC",X"7D",X"F5",X"6D",X"D8",X"7C",
		X"C9",X"7D",X"C4",X"6D",X"F8",X"49",X"B5",X"4D",X"FD",X"E4",X"69",X"FC",X"6D",X"C9",X"49",X"F8",
		X"4D",X"FD",X"DF",X"6D",X"C5",X"4D",X"CD",X"7D",X"E0",X"4D",X"F8",X"49",X"B5",X"6D",X"FD",X"ED",
		X"4D",X"C8",X"75",X"CD",X"7D",X"FE",X"4D",X"C8",X"75",X"CD",X"7D",X"D3",X"6D",X"DC",X"7D",X"F1",
		X"4D",X"CD",X"7F",X"FD",X"CD",X"7D",X"C8",X"75",X"CD",X"7D",X"C8",X"6D",X"F4",X"4D",X"F8",X"49",
		X"CD",X"6D",X"C8",X"75",X"CD",X"7D",X"D0",X"4D",X"E1",X"6D",X"F8",X"69",X"B5",X"4D",X"FD",X"FF",
		X"6D",X"CD",X"7D",X"FF",X"4D",X"C8",X"75",X"CD",X"7D",X"ED",X"4D",X"F8",X"69",X"E5",X"6D",X"E5",
		X"4D",X"F8",X"49",X"B5",X"6D",X"FD",X"CD",X"4D",X"E0",X"6D",X"CD",X"7D",X"CD",X"4D",X"C8",X"75",
		X"CD",X"7D",X"D1",X"4D",X"B5",X"75",X"FD",X"D8",X"7D",X"DC",X"4D",X"C8",X"75",X"D8",X"7D",X"E8",
		X"6D",X"DD",X"7F",X"E9",X"6D",X"E9",X"4D",X"ED",X"5F",X"F8",X"4D",X"E6",X"6D",X"B5",X"4D",X"FD",
		X"F9",X"7D",X"E8",X"6D",X"F5",X"4D",X"F9",X"7D",X"ED",X"6D",X"F8",X"4D",X"F9",X"7D",X"B5",X"6D",
		X"FD",X"8F",X"62",X"99",X"97",X"74",X"C6",X"5C",X"9C",X"FF",X"A2",X"3F",X"B5",X"69",X"F6",X"68",
		X"F6",X"DA",X"DA",X"79",X"A3",X"8F",X"62",X"9D",X"5C",X"78",X"9B",X"1C",X"8A",X"55",X"31",X"09",
		X"29",X"04",X"10",X"77",X"10",X"1D",X"25",X"29",X"05",X"1C",X"77",X"15",X"24",X"77",X"76",X"76",
		X"76",X"76",X"76",X"77",X"34",X"09",X"1D",X"29",X"24",X"10",X"8A",X"8A",X"71",X"B9",X"EF",X"E2",
		X"B6",X"71",X"B9",X"B8",X"E2",X"F3",X"71",X"B9",X"A0",X"E2",X"86",X"73",X"B9",X"0A",X"E2",X"8A",
		X"71",X"B9",X"11",X"E2",X"B6",X"71",X"B9",X"DB",X"C2",X"B6",X"71",X"B9",X"AA",X"C2",X"B5",X"71",
		X"B9",X"B8",X"C2",X"40",X"10",X"1D",X"25",X"29",X"05",X"1C",X"43",X"10",X"77",X"00",X"15",X"24",
		X"11",X"3D",X"1D",X"29",X"01",X"8A",X"AA",X"24",X"3D",X"05",X"77",X"00",X"1D",X"24",X"11",X"3D",
		X"43",X"10",X"77",X"3D",X"09",X"04",X"10",X"05",X"8A",X"8A",X"6B",X"6B",X"6B",X"77",X"00",X"3D",
		X"1D",X"2D",X"05",X"77",X"10",X"3D",X"05",X"43",X"10",X"8A",X"AA",X"77",X"01",X"09",X"29",X"05",
		X"77",X"24",X"09",X"77",X"24",X"3D",X"05",X"8A",X"AA",X"77",X"00",X"1D",X"24",X"11",X"3D",X"05",
		X"10",X"43",X"77",X"31",X"15",X"2D",X"2D",X"6B",X"8A",X"8A",X"3D",X"05",X"2D",X"34",X"77",X"10",
		X"1D",X"25",X"29",X"05",X"1C",X"77",X"34",X"04",X"29",X"11",X"3D",X"8A",X"AA",X"09",X"04",X"24",
		X"77",X"15",X"2D",X"2D",X"77",X"09",X"21",X"77",X"24",X"3D",X"05",X"8A",X"AA",X"01",X"09",X"31",
		X"2D",X"1D",X"29",X"43",X"10",X"77",X"6B",X"6B",X"6B",X"8A",X"8A",X"31",X"05",X"21",X"09",X"30",
		X"05",X"77",X"24",X"3D",X"05",X"1C",X"8A",X"AA",X"25",X"05",X"10",X"24",X"30",X"09",X"1C",X"77",
		X"24",X"3D",X"05",X"8A",X"AA",X"21",X"04",X"30",X"29",X"1D",X"10",X"3D",X"1D",X"29",X"01",X"10",
		X"6B",X"8A",X"8A",X"31",X"05",X"00",X"15",X"30",X"05",X"77",X"09",X"21",X"77",X"05",X"05",X"30",
		X"1D",X"05",X"8A",X"AA",X"10",X"34",X"1D",X"25",X"05",X"30",X"10",X"6B",X"77",X"77",X"77",X"24",
		X"3D",X"05",X"1C",X"8A",X"AA",X"15",X"30",X"05",X"77",X"20",X"05",X"30",X"1C",X"77",X"25",X"05",
		X"15",X"25",X"2D",X"1C",X"57",X"8A",X"8A",X"34",X"04",X"29",X"11",X"3D",X"77",X"09",X"04",X"24",
		X"77",X"31",X"15",X"24",X"10",X"8A",X"AA",X"21",X"09",X"30",X"77",X"31",X"09",X"29",X"04",X"10",
		X"77",X"34",X"09",X"1D",X"29",X"24",X"10",X"6B",X"8A",X"8A",X"31",X"04",X"24",X"77",X"00",X"15",
		X"24",X"11",X"3D",X"77",X"09",X"04",X"24",X"6B",X"8A",X"AA",X"24",X"3D",X"05",X"1C",X"77",X"11",
		X"15",X"29",X"77",X"19",X"1D",X"2D",X"2D",X"57",X"8A",X"8A",X"34",X"04",X"29",X"11",X"3D",X"77",
		X"00",X"1D",X"24",X"11",X"3D",X"77",X"24",X"09",X"8A",X"AA",X"10",X"2D",X"09",X"00",X"77",X"3D",
		X"05",X"30",X"77",X"30",X"05",X"2D",X"05",X"29",X"24",X"4F",X"8A",X"AA",X"2D",X"05",X"10",X"10",
		X"77",X"34",X"04",X"30",X"10",X"04",X"1D",X"24",X"6B",X"8A",X"8A",X"AA",X"47",X"FC",X"F8",X"8B",
		X"FB",X"BF",X"4D",X"AA",X"03",X"FC",X"9E",X"AB",X"03",X"FC",X"1D",X"4C",X"99",X"47",X"FC",X"A4",
		X"60",X"B7",X"39",X"48",X"FB",X"84",X"60",X"AF",X"39",X"48",X"FB",X"97",X"BE",X"E8",X"96",X"E4",
		X"69",X"C2",X"C9",X"5C",X"79",X"9E",X"5C",X"48",X"FB",X"15",X"0C",X"45",X"55",X"4D",X"8F",X"6B",
		X"F8",X"53",X"62",X"AE",X"9B",X"C7",X"B6",X"EA",X"8F",X"6F",X"F8",X"53",X"E7",X"18",X"F9",X"AE",
		X"BB",X"E2",X"DF",X"A3",X"BF",X"FC",X"AA",X"A6",X"FC",X"F0",X"8B",X"F1",X"8B",X"55",X"F0",X"8B",
		X"F1",X"8B",X"A2",X"BF",X"FC",X"4B",X"E0",X"AF",X"FB",X"8B",X"AB",X"A6",X"FC",X"E2",X"DF",X"A3",
		X"6B",X"F8",X"0D",X"5C",X"9C",X"FF",X"0D",X"15",X"05",X"1C",X"97",X"F1",X"BB",X"8F",X"80",X"C2",
		X"9F",X"DA",X"40",X"10",X"C8",X"19",X"51",X"C9",X"19",X"73",X"DB",X"BF",X"98",X"D6",X"30",X"77");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
